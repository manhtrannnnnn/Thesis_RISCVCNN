`timescale 1 ns / 1 ps

`define TIME_TO_REPEAT 6
// `define FCL_TC0
`define ML_TC1
// `define CL_TC2
     
module al_accel_tb;
    localparam 
        CONV    = 4'd 0,
        DENSE   = 4'd 1,
        MIXED   = 4'd 2;

    localparam 
        RELU    = 4'd0,
        RELU6   = 4'd1,
        SIGMOID = 4'd2,
        TANH    = 4'd3,
        NO_FUNC = 4'd4;

    // Mandatory Sigs Control
    reg clk;
	always #5 clk = (clk === 1'b0); 

    reg resetn;
    initial begin
        resetn = 1'b 0;
        #42
        resetn = 1'b 1;
    end

    // SoC Ctrl Sigs
    reg  [31:0] al_accel_cfgreg_di;
    reg  [ 4:0] al_accel_cfgreg_sel;
    reg         al_accel_cfgreg_wenb;
    reg         al_accel_flow_enb;
    reg         al_accel_mem_read_ready;
    reg         al_accel_mem_write_ready;

    wire [31:0] al_accel_raddr, al_accel_waddr;
    wire        al_accel_renb , al_accel_wenb;
    wire [ 3:0] al_accel_wstrb;
    wire [31:0] al_accel_rdata, al_accel_wdata;
    wire al_accel_cal_fin;

// Convolutional Layer
`ifdef CL_TC0
/* Test case 0 */
     /* 
        Description:
           - Input Feature Map's size : 13 x 13 x 32     => 5048 -> 1352
           - Kernel's size            : 3 x 3 x 32 x 32 => 9216 -> 2304
           - Output Feature Map's size: 11 x 11 x 32     => 3872 -> 968
           - Bias's size              : 32 x 1         =>  32
           - Partial-Sum's size       : 6 x 6 x 6 x 4 => 864
    */

    localparam 
        IFM_SIZE = 13 * 13 * 32     + 1,
        KER_SIZE = 3 * 3 * 32 * 32 + 2,
        OFM_SIZE = 11 * 11 * 32     + 2,
        BIS_SIZE = 32,
        PAS_SIZE = 5 * 5 * 6;

    initial begin
        // al_accel_mem_read_ready = 1'b 0;
        // al_accel_mem_write_ready = 1'b 0;
        // #10
        // repeat (2000) @(posedge clk) begin
        //     #2 al_accel_mem_read_ready = $random;
        // end
        // #10 
        al_accel_mem_read_ready    = 1'b 1;
        al_accel_mem_write_ready   = 1'b 1;
    end

    initial begin
        al_accel_cfgreg_di   = 32'd 0; al_accel_cfgreg_sel = 5'd 0; 
        al_accel_cfgreg_wenb =  1'd 0;
        al_accel_flow_enb    =  1'b 0;
        #42
        al_accel_cfgreg_wenb =  1'd 1;
    // Config Data
        #10 // i_base_addr
        al_accel_cfgreg_di   = 32'd 0;       al_accel_cfgreg_sel = 5'd 0; 

        #10 // kw_base_addr
        al_accel_cfgreg_di   = 32'd 6000;       al_accel_cfgreg_sel = 5'd 1; 

        #10 // o_base_addr
        al_accel_cfgreg_di   = 32'd 16000;       al_accel_cfgreg_sel = 5'd 2; 

        #10 // b_base_addr
        al_accel_cfgreg_di   = 32'd 5600;       al_accel_cfgreg_sel = 5'd 3; 

        #10 // ps_base_addr
        al_accel_cfgreg_di   = 32'd 20000;       al_accel_cfgreg_sel = 5'd 4; 

        #10 // {stride_height, stride_width, cfg_act_func_typ, cfg_layer_typ}
        al_accel_cfgreg_di   = {16'd 0, 4'd 1, 4'd 1, RELU, CONV}; al_accel_cfgreg_sel = 5'd 5; 

        #10 // {weight_kernel_patch_height, weight_kernel_patch_width}
        al_accel_cfgreg_di   = {16'd 3, 16'd 3}; al_accel_cfgreg_sel = 5'd 6; 

        #10 // {nok_ofm_depth, kernel_ifm_depth} 
        al_accel_cfgreg_di   = {16'd 6, 16'd 3}; al_accel_cfgreg_sel = 5'd 7;
        
        #10 // {ifm_height, ifm_width}  
        al_accel_cfgreg_di   = {16'd 7, 16'd 7}; al_accel_cfgreg_sel = 5'd 8;

        #10 // {ofm_height, ofm_width}
        al_accel_cfgreg_di   = {16'd 5, 16'd 5}; al_accel_cfgreg_sel = 5'd 9;

        #10 // {output2D_size, input2D_size}  
        al_accel_cfgreg_di   = {16'd 25, 16'd 49}; al_accel_cfgreg_sel = 5'd 10;

        #10 // kernel3D_size
        al_accel_cfgreg_di   = {16'd  0, 16'd 27}; al_accel_cfgreg_sel = 5'd 11;

    // Output Quantize Buffer
        #10 // output_quant_sel 0
        al_accel_cfgreg_di   = {24'd 0, 8'd 0} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1689551407 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 1
        al_accel_cfgreg_di   = {24'd 0, 8'd 1} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1204010513 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 2
        al_accel_cfgreg_di   = {24'd 0, 8'd 2} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2140008272 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 3
        al_accel_cfgreg_di   = {24'd 0, 8'd 3} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1909323516 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 4
        al_accel_cfgreg_di   = {24'd 0, 8'd 4} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1725018846 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 5
        al_accel_cfgreg_di   = {24'd 0, 8'd 5} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2048260720 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 6
        al_accel_cfgreg_di   = {24'd 0, 8'd 6} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2126767021 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 7
        al_accel_cfgreg_di   = {24'd 0, 8'd 7} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1808926684 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 8
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1463903110 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 9
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1253391477 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 10
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1548369488 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 11
        al_accel_cfgreg_di   = {24'd 0, 8'd 11} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1854827854 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 12
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1089899269 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 13
        al_accel_cfgreg_di   = {24'd 0, 8'd 13} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1700026496 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 14
        al_accel_cfgreg_di   = {24'd 0, 8'd 14} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2095039993 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 15
        al_accel_cfgreg_di   = {24'd 0, 8'd 15} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1336030234 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 16
        al_accel_cfgreg_di   = {24'd 0, 8'd 16} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1663159508 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 17
        al_accel_cfgreg_di   = {24'd 0, 8'd 17} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1997878220 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 18
        al_accel_cfgreg_di   = {24'd 0, 8'd 18} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1660705979 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 19
        al_accel_cfgreg_di   = {24'd 0, 8'd 19} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1740647325 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 20
        al_accel_cfgreg_di   = {24'd 0, 8'd 20} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1385151967 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 21
        al_accel_cfgreg_di   = {24'd 0, 8'd 21} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1207776079 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 22
        al_accel_cfgreg_di   = {24'd 0, 8'd 22} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1712031603 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 23
        al_accel_cfgreg_di   = {24'd 0, 8'd 23} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1593821800 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 24
        al_accel_cfgreg_di   = {24'd 0, 8'd 24} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1368997244 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 25
        al_accel_cfgreg_di   = {24'd 0, 8'd 25} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1466326579 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 26
        al_accel_cfgreg_di   = {24'd 0, 8'd 26} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1582443027 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 27
        al_accel_cfgreg_di   = {24'd 0, 8'd 27} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1558951275 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 28
        al_accel_cfgreg_di   = {24'd 0, 8'd 28} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1682677520 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 29
        al_accel_cfgreg_di   = {24'd 0, 8'd 29} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1747796433 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 30
        al_accel_cfgreg_di   = {24'd 0, 8'd 30} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1716120888 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 31
        al_accel_cfgreg_di   = {24'd 0, 8'd 31} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1544083328 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

    // Data Offset
        #10 // input_offset
        al_accel_cfgreg_di   = 32'd 0; al_accel_cfgreg_sel = 5'd 15;
        #10 // output_offset
        al_accel_cfgreg_di   = 32'd 0; al_accel_cfgreg_sel = 5'd 16;

    // Flow Run
        #10
        al_accel_cfgreg_wenb =  1'd 0;
        #10 
        al_accel_flow_enb    =  1'd 1;
        // #1000
        // al_accel_flow_enb    =  1'd 0;
        // #200
        al_accel_flow_enb    =  1'd 1;
		// repeat (2000) @(posedge clk) begin
        //     #2 al_accel_flow_enb = $random;
        // end
        // #10 
        al_accel_flow_enb    =  1'd 1;
    end

    reg [IFM_SIZE     * 8 - 1:0] input_data ; // Size: 7 x 7 x 3
    reg [KER_SIZE * 8 - 1:0] filter_data; // Size: 3 x 3 x 3 x 6
    reg [BIS_SIZE * 32                 - 1:0] bias_data  ; // Size: 6
    integer i;
    initial begin
        for (i = 0; i < 8192; i = i + 1)
            ram.mem[i] = 32'd 0;

        // Input Initilization
        input_data = {
             -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd90, -8'd46, -8'd63, -8'd110, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd27, 8'd58, 8'd42, 8'd63, 8'd63, 8'd69, 8'd65, 8'd61, -8'd23, -8'd128, -8'd128, -8'd128, -8'd128, -8'd127, -8'd128, -8'd128, -8'd111, -8'd93, -8'd81, -8'd73, -8'd13, -8'd43, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd110, -8'd3, -8'd34, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd41, -8'd11, -8'd96, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd111, -8'd26, -8'd46, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd126, -8'd20, 8'd4, -8'd103, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd66, 8'd9, -8'd36, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd108, 8'd11, -8'd24, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd44, 8'd3, -8'd52, -8'd119, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd56, -8'd35, -8'd117, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd98, -8'd102, -8'd119, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd40, -8'd2, -8'd5, -8'd21, -8'd39, -8'd39, -8'd39, -8'd40, -8'd114, -8'd128, -8'd128, -8'd128, -8'd128, -8'd70, -8'd36, -8'd15, 8'd1, -8'd2, -8'd1, 8'd23, 8'd27, -8'd65, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd120, -8'd115, -8'd107, -8'd10, -8'd17, -8'd82, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd52, -8'd11, -8'd28, -8'd119, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd108, -8'd20, -8'd15, -8'd89, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd126, -8'd50, -8'd14, -8'd44, -8'd123, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd73, -8'd14, -8'd16, -8'd93, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd106, -8'd13, -8'd15, -8'd59, -8'd126, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd52, 8'd28, -8'd14, -8'd115, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd28, 8'd13, -8'd32, -8'd122, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd97, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd84, -8'd99, -8'd99, -8'd99, -8'd99, -8'd111, -8'd94, -8'd110, -8'd89, -8'd92, -8'd91, -8'd94, -8'd115, -8'd6, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd96, -8'd97, -8'd95, -8'd128, -8'd11, -8'd10, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd109, -8'd128, -8'd6, -8'd75, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd128, 8'd0, -8'd15, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd112, -8'd119, -8'd1, -8'd87, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd128, -8'd8, -8'd22, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd128, -8'd24, -8'd8, -8'd92, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd110, -8'd128, -8'd11, -8'd65, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99, -8'd128, -8'd57, -8'd15, -8'd82, -8'd99, -8'd99, -8'd99, -8'd99, -8'd99,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd117, -8'd109, -8'd119, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd75, -8'd2, -8'd27, -8'd50, -8'd59, -8'd58, -8'd55, -8'd57, -8'd59, -8'd128, -8'd128, -8'd128, -8'd128, -8'd64, -8'd25, -8'd12, 8'd4, 8'd3, 8'd8, 8'd11, 8'd36, -8'd19, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd120, -8'd114, -8'd110, -8'd55, 8'd26, -8'd56, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd121, 8'd37, 8'd23, -8'd117, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd47, 8'd25, -8'd68, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd114, 8'd29, 8'd7, -8'd125, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd25, 8'd34, -8'd77, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd60, 8'd41, -8'd25, -8'd127, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd121, 8'd26, 8'd26, -8'd105, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd59, 8'd59, 8'd11, -8'd120, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd71, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd70, -8'd128, -8'd128, -8'd127, -8'd113, -8'd113, -8'd113, -8'd115, -8'd89, -8'd78, -8'd78, -8'd78, -8'd78, -8'd94, -8'd97, -8'd118, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd89, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd73, -8'd74, -8'd128, -8'd75, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd73, -8'd128, -8'd78, -8'd76, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd73, -8'd85, -8'd128, -8'd76, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd77, -8'd70, -8'd128, -8'd77, -8'd75, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd69, -8'd95, -8'd126, -8'd75, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd73, -8'd70, -8'd128, -8'd74, -8'd76, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd74, -8'd128, -8'd128, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78, -8'd89, -8'd128, -8'd71, -8'd76, -8'd78, -8'd78, -8'd78, -8'd78, -8'd78,, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd97, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd93, -8'd90, -8'd90, -8'd90, -8'd90, -8'd107, -8'd102, -8'd126, -8'd128, -8'd127, -8'd128, -8'd128, -8'd128, -8'd60, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd99, -8'd93, -8'd49, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd128, -8'd44, -8'd72, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd117, -8'd70, -8'd43, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd91, -8'd128, -8'd43, -8'd78, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd128, -8'd58, -8'd44, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd102, -8'd120, -8'd45, -8'd83, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd128, -8'd66, -8'd68, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90, -8'd114, -8'd128, -8'd46, -8'd79, -8'd90, -8'd90, -8'd90, -8'd90, -8'd90,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd67, -8'd30, -8'd60, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd119, -8'd113, -8'd113, -8'd113, -8'd113, -8'd33, 8'd9, 8'd24, 8'd19, 8'd7, 8'd1, 8'd6, -8'd56, -8'd59, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd111, -8'd100, -8'd93, -8'd88, -8'd128, -8'd38, -8'd61, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd123, -8'd51, -8'd29, -8'd100, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd128, -8'd39, -8'd68, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd126, -8'd54, -8'd44, -8'd107, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd89, -8'd27, -8'd70, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd128, -8'd25, -8'd32, -8'd109, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd124, -8'd92, -8'd76, -8'd102, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113, -8'd30, 8'd29, -8'd17, -8'd104, -8'd113, -8'd113, -8'd113, -8'd113, -8'd113,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd95, -8'd88, -8'd104, -8'd124, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd11, 8'd16, 8'd12, -8'd6, -8'd18, -8'd17, -8'd19, -8'd21, -8'd108, -8'd128, -8'd128, -8'd128, -8'd128, -8'd43, -8'd18, 8'd10, 8'd24, 8'd17, 8'd18, 8'd38, 8'd74, -8'd64, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd127, -8'd114, -8'd109, -8'd102, 8'd31, 8'd36, -8'd89, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd32, 8'd34, -8'd8, -8'd123, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd108, 8'd26, 8'd31, -8'd99, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd125, -8'd24, 8'd30, -8'd29, -8'd123, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd61, 8'd30, 8'd23, -8'd102, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd104, 8'd24, 8'd40, -8'd57, -8'd125, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd33, 8'd70, 8'd16, -8'd118, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd1, 8'd58, -8'd17, -8'd125, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd93, -8'd81, -8'd99, -8'd123, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd6, 8'd46, 8'd45, 8'd24, 8'd7, 8'd6, 8'd3, 8'd2, -8'd96, -8'd128, -8'd128, -8'd128, -8'd128, -8'd28, 8'd1, 8'd34, 8'd51, 8'd53, 8'd53, 8'd59, 8'd108, -8'd56, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd126, -8'd111, -8'd106, -8'd101, 8'd57, 8'd71, -8'd79, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd17, 8'd74, 8'd9, -8'd120, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd113, 8'd56, 8'd71, -8'd91, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd126, 8'd0, 8'd59, -8'd13, -8'd124, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd59, 8'd72, 8'd63, -8'd94, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd108, 8'd47, 8'd72, -8'd41, -8'd125, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd20, 8'd109, 8'd53, -8'd119, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd15, 8'd99, -8'd2, -8'd123, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd40, 8'd18, -8'd11, -8'd80, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd18, 8'd14, 8'd46, 8'd52, 8'd42, 8'd42, 8'd42, 8'd36, -8'd38, -8'd104, -8'd104, -8'd104, -8'd104, -8'd118, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd96, -8'd95, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd77, -8'd51, -8'd120, -8'd106, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd47, -8'd61, -8'd128, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd77, -8'd57, -8'd128, -8'd105, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd100, -8'd39, -8'd52, -8'd125, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd57, -8'd27, -8'd128, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd77, -8'd42, -8'd108, -8'd110, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd50, -8'd62, -8'd106, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd99, -8'd128, -8'd128, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd104, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd112, -8'd68, -8'd78, -8'd113, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd35, 8'd19, 8'd9, 8'd16, 8'd15, 8'd18, 8'd17, 8'd10, -8'd45, -8'd128, -8'd128, -8'd128, -8'd128, -8'd57, -8'd39, -8'd17, 8'd2, 8'd7, 8'd17, 8'd12, 8'd56, -8'd22, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd127, -8'd119, -8'd114, -8'd113, 8'd26, 8'd63, -8'd77, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd60, 8'd71, 8'd25, -8'd124, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd124, 8'd25, 8'd59, -8'd91, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd43, 8'd59, 8'd6, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd93, 8'd73, 8'd67, -8'd98, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd121, 8'd20, 8'd68, -8'd43, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd61, 8'd91, 8'd56, -8'd113, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd35, 8'd78, 8'd5, -8'd125, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd93, -8'd84, -8'd103, -8'd125, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd31, 8'd2, 8'd10, 8'd6, -8'd4, -8'd5, -8'd8, -8'd9, -8'd94, -8'd128, -8'd128, -8'd128, -8'd128, -8'd72, -8'd48, -8'd25, -8'd8, 8'd1, 8'd3, 8'd17, 8'd46, -8'd75, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd127, -8'd121, -8'd118, -8'd109, 8'd18, 8'd5, -8'd93, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd26, 8'd18, -8'd47, -8'd121, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd111, 8'd9, 8'd6, -8'd97, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd126, -8'd13, 8'd13, -8'd61, -8'd126, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd59, 8'd16, 8'd2, -8'd100, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd107, 8'd17, 8'd9, -8'd76, -8'd127, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd28, 8'd50, -8'd9, -8'd119, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd8, 8'd35, -8'd56, -8'd122, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd108, -8'd91, -8'd100, -8'd122, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd28, -8'd2, -8'd9, -8'd11, -8'd19, -8'd19, -8'd20, -8'd21, -8'd87, -8'd128, -8'd128, -8'd128, -8'd128, -8'd63, -8'd47, -8'd25, -8'd4, -8'd1, 8'd1, -8'd5, 8'd35, -8'd67, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd126, -8'd119, -8'd116, -8'd114, 8'd21, 8'd27, -8'd102, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd51, 8'd31, -8'd31, -8'd124, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd123, 8'd16, 8'd27, -8'd108, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd34, 8'd25, -8'd49, -8'd127, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd94, 8'd32, 8'd23, -8'd111, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd121, 8'd18, 8'd28, -8'd80, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd53, 8'd47, 8'd10, -8'd122, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd24, 8'd37, -8'd46, -8'd125, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd115, -8'd104, -8'd127, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd49, -8'd58, -8'd80, -8'd69, -8'd59, -8'd55, -8'd51, -8'd59, -8'd84, -8'd128, -8'd128, -8'd128, -8'd128, -8'd96, -8'd128, -8'd128, -8'd128, -8'd128, -8'd122, -8'd120, -8'd105, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd8, 8'd5, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd99, 8'd12, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd9, -8'd17, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd77, 8'd11, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd4, -8'd29, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd8, 8'd17, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd101, -8'd19, -8'd115, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd55, -8'd45, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd112, -8'd72, -8'd81, -8'd116, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd30, 8'd12, -8'd1, 8'd10, 8'd10, 8'd14, 8'd12, 8'd7, -8'd52, -8'd128, -8'd128, -8'd128, -8'd128, -8'd50, -8'd46, -8'd24, -8'd7, -8'd1, 8'd10, 8'd6, 8'd40, -8'd41, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd120, -8'd114, -8'd116, 8'd34, 8'd65, -8'd95, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd51, 8'd73, 8'd3, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd125, 8'd33, 8'd59, -8'd108, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd34, 8'd60, -8'd14, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd89, 8'd75, 8'd64, -8'd114, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd122, 8'd29, 8'd68, -8'd62, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd53, 8'd88, 8'd39, -8'd122, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd23, 8'd67, -8'd18, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd44, -8'd66, -8'd91, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd107, -8'd94, -8'd94, -8'd94, -8'd94, -8'd22, 8'd21, 8'd33, 8'd15, 8'd17, 8'd16, 8'd7, -8'd71, -8'd79, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd91, -8'd82, -8'd69, -8'd66, -8'd79, -8'd124, -8'd69, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd86, -8'd120, -8'd51, -8'd81, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd75, -8'd98, -8'd62, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd98, -8'd128, -8'd63, -8'd83, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd81, -8'd119, -8'd71, -8'd64, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd103, -8'd119, -8'd55, -8'd87, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd83, -8'd120, -8'd128, -8'd88, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd6, 8'd2, -8'd40, -8'd86, -8'd94, -8'd94, -8'd94, -8'd94, -8'd94, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd93, -8'd59, -8'd72, -8'd115, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd43, 8'd18, 8'd17, 8'd25, 8'd23, 8'd26, 8'd22, 8'd23, -8'd50, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd89, -8'd87, -8'd79, -8'd79, 8'd20, -8'd28, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd118, -8'd53, -8'd30, -8'd93, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd97, -8'd47, -8'd39, -8'd122, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd118, -8'd66, -8'd42, -8'd99, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd127, -8'd72, -8'd43, -8'd48, -8'd126, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd104, -8'd40, -8'd45, -8'd104, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd117, -8'd52, -8'd39, -8'd85, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd100, -8'd20, 8'd11, -8'd115, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd115, -8'd43, -8'd50, -8'd124, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd80, -8'd40, -8'd63, -8'd111, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd18, 8'd51, 8'd42, 8'd47, 8'd56, 8'd61, 8'd56, 8'd54, -8'd43, -8'd128, -8'd128, -8'd128, -8'd128, -8'd118, -8'd128, -8'd128, -8'd106, -8'd89, -8'd77, -8'd59, -8'd16, -8'd63, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd103, 8'd29, -8'd4, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd29, 8'd18, -8'd91, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd104, 8'd5, -8'd22, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd125, -8'd8, 8'd30, -8'd101, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd59, 8'd38, -8'd22, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd102, 8'd39, 8'd9, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd31, 8'd35, -8'd44, -8'd126, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd28, -8'd3, -8'd114, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd98, -8'd91, -8'd106, -8'd122, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd70, -8'd21, -8'd13, -8'd20, -8'd29, -8'd29, -8'd29, -8'd32, -8'd90, -8'd126, -8'd126, -8'd126, -8'd126, -8'd104, -8'd64, -8'd50, -8'd34, -8'd29, -8'd27, -8'd5, -8'd3, -8'd52, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd122, -8'd117, -8'd106, -8'd43, -8'd39, -8'd69, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd66, -8'd42, -8'd37, -8'd113, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd107, -8'd53, -8'd41, -8'd75, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd123, -8'd63, -8'd42, -8'd47, -8'd120, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd75, -8'd37, -8'd38, -8'd80, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd105, -8'd42, -8'd34, -8'd56, -8'd122, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd66, 8'd3, -8'd26, -8'd105, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126, -8'd59, -8'd16, -8'd39, -8'd116, -8'd126, -8'd126, -8'd126, -8'd126, -8'd126,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd109, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd31, -8'd79, -8'd82, -8'd125, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd58, -8'd61, -8'd43, -8'd38, -8'd57, -8'd68, -8'd16, -8'd2, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd126, -8'd123, -8'd113, -8'd42, -8'd78, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd53, -8'd49, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd115, -8'd29, -8'd87, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd59, -8'd60, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd69, -8'd36, -8'd122, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd111, -8'd52, -8'd62, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd53, -8'd35, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd23, -8'd34, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd77, -8'd98, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd109, -8'd101, -8'd101, -8'd101, -8'd101, 8'd7, 8'd43, 8'd47, 8'd48, 8'd54, 8'd49, 8'd31, -8'd57, -8'd98, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd97, -8'd79, -8'd67, -8'd58, -8'd109, -8'd80, -8'd80, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd109, -8'd98, -8'd59, -8'd93, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd120, -8'd79, -8'd77, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd112, -8'd105, -8'd79, -8'd91, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd102, -8'd128, -8'd66, -8'd77, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd128, -8'd71, -8'd58, -8'd95, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd110, -8'd128, -8'd124, -8'd97, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101, -8'd19, 8'd13, -8'd31, -8'd94, -8'd101, -8'd101, -8'd101, -8'd101, -8'd101,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd117, -8'd126, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd102, -8'd123, -8'd121, -8'd128, -8'd128, -8'd128, -8'd78, -8'd45, -8'd128, -8'd128, -8'd128, -8'd128, -8'd127, -8'd79, -8'd101, -8'd77, -8'd93, -8'd79, -8'd73, 8'd18, 8'd7, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd126, -8'd128, -8'd125, -8'd128, 8'd42, -8'd46, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd25, 8'd39, -8'd127, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd44, -8'd65, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd28, 8'd39, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd58, 8'd36, -8'd77, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd38, -8'd2, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd88, 8'd33, -8'd112, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd14, 8'd29, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,  -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd122, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd16, 8'd3, -8'd9, -8'd61, -8'd87, -8'd91, -8'd87, -8'd94, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd44, -8'd23, 8'd10, 8'd21, 8'd22, 8'd17, 8'd34, 8'd6, -8'd109, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd125, -8'd116, -8'd114, -8'd113, -8'd35, -8'd57, -8'd102, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd42, -8'd31, -8'd82, -8'd120, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd117, -8'd23, -8'd51, -8'd104, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd127, -8'd55, -8'd47, -8'd100, -8'd127, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd64, -8'd33, -8'd51, -8'd104, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd111, -8'd35, -8'd50, -8'd87, -8'd127, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd41, -8'd15, -8'd96, -8'd126, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd10, 8'd12, -8'd77, -8'd121, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128
        };
        for (i = 0; i < (13 * 13 * 32 + 1); i = i + 4) begin
            ram.mem[0 + (i / 4)][ 7: 0] = input_data[8*((7 * 7 * 3 + 1) - 1 - i) +: 8];
            ram.mem[0 + (i / 4)][15: 8] = input_data[8*((7 * 7 * 3 + 1) - 2 - i) +: 8];
            ram.mem[0 + (i / 4)][23:16] = input_data[8*((7 * 7 * 3 + 1) - 3 - i) +: 8];
            ram.mem[0 + (i / 4)][31:24] = input_data[8*((7 * 7 * 3 + 1) - 4 - i) +: 8];
        end

        // Kernel 
        filter_data = {
        -79, -97, -56, -108, -102, 2, -70, 60, -66, 
        -123, -100, -71, 84, -83, -36, 3, -116, 34, 
        38, -87, 57, 60, 21, -3, -49, -82, -57, 
        65, 89, -62, -126, -87, -25, -127, -62, 73, 
        -32, 64, 48, -10, 7, 32, -54, -80, 92, 
        4, 33, -65, 87, 2, -73, -107, -15, -77, 
        40, 87, -29, -106, -70, -19, -4, 64, -118, 
        79, -64, 82, -40, 78, 0, -29, 95, -94, 
        7, 23, -57, -118, -90, 36, -115, 15, -58, 
        -8, -74, 7, -104, -34, -36, -113, 90, -96, 
        -73, -17, 44, 107, -87, -38, -93, 93, 2, 
        -121, 37, 68, -62, 3, -113, 84, -57, -86, 
        54, -92, -40, -109, 50, 16, 87, 64, 41, 
        71, 32, 2, -24, -55, -101, 85, -52, 88, 
        -6, 34, -83, 55, -58, -14, -5, 70, -118, 
        -18, 14, 8, 8, 30, -99, 83, -2, -42, 
        75, -25, -41, 4, -3, -79, 40, -104, -24, 
        -70, 92, 52, -74, 13, 99, -73, -73, 19, 
        -28, -32, -71, -4, -4, 77, 7, 54, -46, 
        81, -65, 15, -68, 1, 44, 91, 84, 7, 
        24, -92, -78, 17, -109, -69, -74, -49, 57, 
        -29, 12, -28, -92, 44, -119, 39, 20, 43, 
        -101, 70, 63, -7, 39, 81, -104, -46, -11, 
        62, 98, 54, 61, -56, -75, 84, 82, 41, 
        -68, -66, 48, -119, -120, -46, -52, -47, -118, 
        31, 33, 102, 81, 27, -96, -15, 39, 61, 
        -23, 33, 75, 106, -68, -46, -4, 25, -9, 
        -63, -32, -14, 97, -15, -109, -33, -100, 101, 
        -71, 10, 82, -71, 51, 110, -25, 13, -21, 
        29, 8, 71, -3, 36, -38, -67, -58, -42, 
        73, 68, 31, -108, -107, -102, -64, -88, 69, 
        12, 88, -30, 95, -115, 30, 14, -20, 53, 
        45, -17, -48, 23, -8, -35, -33, -106, -15, 
        41, 3, 9, 20, 11, -7, -2, -47, -2, 
        27, 4, 1, 20, 32, 13, 18, 20, 21, 
        24, 31, -5, 29, 5, -27, 25, 0, -20, 
        21, -13, 13, -6, -14, 1, 19, 10, -16, 
        -13, 8, 20, -8, 14, 10, 14, 26, 17, 
        3, -13, 16, 22, 30, -4, 11, 19, -14, 
        -8, 13, -17, 15, 19, -12, 6, 13, -2, 
        25, 0, 7, 20, 5, -1, 21, -3, 8, 
        29, 27, 10, 45, -9, -16, -27, -52, -17, 
        -19, -14, -13, 2, -3, -10, 18, 9, -3, 
        39, 17, -3, 26, 7, -50, 11, -52, 18, 
        -47, -51, -60, -53, -22, -10, -47, -47, -26, 
        14, -8, -6, 5, 20, 12, 16, 12, 8, 
        39, 35, -18, 26, -19, -45, 5, -57, -18, 
        31, 24, -11, 26, -10, -39, -21, -56, -19, 
        24, 4, -22, 37, -20, -32, -18, -41, -12, 
        19, -60, -127, -41, -62, 14, -70, -43, 57, 
        15, 13, 3, 11, 15, -8, 6, 1, 12, 
        18, -10, 1, -10, 8, -7, 15, 7, -6, 
        52, 34, -13, 22, -16, -7, 19, -65, -24, 
        -18, -14, 5, 8, -9, -18, 10, -11, 18, 
        51, 12, -40, 13, -27, -32, -21, -71, -27, 
        32, 7, -54, -5, -18, -22, -61, -64, 10, 
        33, 25, 17, 30, -3, -8, 14, -25, -15, 
        2, -13, 7, -1, -16, 18, -1, 15, -17, 
        9, 9, -43, -3, -69, -49, -85, -114, 16, 
        -7, -10, -5, 16, -1, -13, -12, 13, 0, 
        3, 16, -19, -13, -6, 0, 17, -11, -11, 
        -64, 3, -1, -15, -10, -24, 22, -9, -10, 
        74, 36, 14, 29, 24, -22, 27, -24, -49, 
        10, -11, -37, 23, -27, -53, -32, -11, 11, 
        6, -7, -3, -20, -36, -3, -25, -22, -17, 
        -37, 15, 6, -16, 12, 39, -23, 14, 41, 
        -7, 0, -30, 6, -5, -2, 12, 16, 2, 
        -11, -30, 1, 7, -35, 23, 8, -27, 19, 
        1, 16, -17, -14, -12, -10, -16, 16, 1, 
        1, 20, -11, 7, 41, -49, -17, 8, -28, 
        31, 30, -49, 3, 4, -29, 29, 21, -20, 
        -14, 13, 14, -5, -1, -20, 14, -1, -5, 
        -10, -45, -6, 7, -42, -21, 16, -28, 4, 
        -35, -8, 43, -33, -3, 36, -43, -29, 47, 
        -22, 16, 22, 6, -8, -21, 5, 17, -7, 
        -24, -7, 55, -27, -2, 29, -45, -13, 73, 
        14, -29, -48, 20, -49, -46, 0, -55, -49, 
        -22, -17, -16, 13, 10, 8, 18, 6, -11, 
        -28, -24, 29, -8, -15, 32, -32, -19, 42, 
        -50, 23, 41, -14, 3, 29, -52, -2, 28, 
        -54, -14, 43, -22, 8, 23, -17, -39, 22, 
        0, -23, 39, -43, 9, -47, -27, -66, -57, 
        18, -17, 17, 4, -16, -4, -4, -10, -8, 
        19, -14, -6, -4, 8, 15, 17, -4, 3, 
        -42, -5, 44, -1, -8, 42, -31, -25, 41, 
        -31, 8, 4, 14, 22, -26, 32, 4, 3, 
        -9, -55, 30, -18, -41, 15, -40, -38, 46, 
        -30, 5, 2, -7, -29, 9, -43, -9, 28, 
        -28, -9, 8, 17, -9, 22, -10, 14, 3, 
        -6, -20, 8, -14, -13, 12, -15, -21, -5, 
        -85, 11, 85, -62, 10, 79, -36, 26, 127, 
        -20, -2, -9, 6, -20, -12, 6, 5, 3, 
        17, -5, 9, 13, 10, 21, -13, -3, 2, 
        -11, -12, -102, 14, -44, -66, 51, 12, -31, 
        14, -46, 71, 12, -61, 37, -1, -111, -8, 
        -44, 13, 17, -33, 4, 32, -12, 12, 38, 
        -16, -50, -14, 45, 10, -71, 24, 51, 4, 
        -1, 12, 53, -20, -40, -50, 60, 32, 7, 
        -24, -18, 13, -58, -27, -1, -10, -10, -35, 
        14, -13, 36, -33, -12, -48, 37, 47, -1, 
        3, -10, -23, -19, -6, 21, 22, 11, 8, 
        25, 19, 27, 37, 18, -15, -24, 12, -9, 
        0, 16, 16, -18, 11, -27, 14, -18, -31, 
        -9, 8, -3, 14, 11, 1, 7, 12, 8, 
        20, 48, 9, -12, -48, -3, 36, -14, -54, 
        -30, -1, 22, -34, -60, -46, 67, 15, -37, 
        20, -18, -19, -6, -13, 9, 3, -8, -24, 
        -35, -1, 47, -58, -85, -63, 43, 58, -18, 
        -13, -15, -59, 98, 62, -10, -8, -3, -7, 
        -11, -8, -5, -1, 17, 19, -23, 23, 18, 
        -1, -19, 39, -5, -30, -36, 57, 16, -23, 
        -29, -6, 22, 3, -38, -59, 34, 15, -33, 
        -46, -25, 18, -35, -37, -60, 37, 40, -12, 
        -39, -127, 21, -71, -91, -61, -21, -52, -68, 
        17, -9, -15, 17, -11, -15, -24, 8, -12, 
        -12, 12, -1, -6, -12, -9, -5, -6, -1, 
        -17, -33, 17, -37, -27, -77, 19, 25, -25, 
        20, 9, 2, -17, 15, 28, 38, -19, -24, 
        -76, -36, -17, 59, -6, -70, 54, 43, 4, 
        -43, -66, 10, 48, -5, -37, 50, 8, -15, 
        17, -8, 17, 11, 14, -21, 59, 22, 32, 
        4, 9, 23, 12, -22, -15, 14, 4, -7, 
        -41, 6, 19, -75, -67, 49, 82, 127, 31, 
        -1, 6, -11, -6, 12, -24, 23, 2, 12, 
        15, -3, 7, 7, 15, -13, -9, -23, -16, 
        102, 42, 8, 15, 44, 44, 35, 20, -28, 
        -80, -72, -16, -36, -42, -91, 12, 38, -40, 
        5, 10, 52, -65, -113, -40, 59, 16, -50, 
        -56, -56, -89, 32, -73, 64, -72, 99, -33, 
        -5, -56, 40, 29, -108, 101, -66, 96, 7, 
        -33, -111, 69, 54, 86, -63, 1, -95, -6, 
        -1, 70, 6, 55, 33, 90, -12, -22, -81, 
        1, 100, -35, -4, 58, -43, -2, 57, -37, 
        -115, 70, 19, 29, -46, -77, -119, -3, -5, 
        34, -46, -4, 10, -99, -53, 81, -7, -18, 
        -105, 33, -81, -32, 62, 78, 16, 52, -100, 
        -58, -99, -93, 36, -59, -59, 78, -92, -64, 
        -47, -94, 53, -50, 4, 0, 65, 1, 1, 
        73, 77, -42, -36, 88, 44, -10, 48, -55, 
        -69, 7, -81, -127, -77, 43, -17, -49, -99, 
        57, 63, -76, 39, -116, 56, -64, -59, -13, 
        -5, 28, 10, 37, 32, 92, 8, 58, -63, 
        -108, -39, 24, -67, -106, -93, 39, 40, -84, 
        51, -23, -24, 74, 22, -111, -95, -83, -73, 
        -48, 29, 19, -4, -99, 78, -119, 51, -64, 
        69, 58, -46, 65, -8, 104, 46, 61, -11, 
        -77, -15, -45, 83, 38, -36, -79, -73, 79, 
        30, -102, -74, 89, 91, -31, 45, 23, -35, 
        41, -38, 80, 2, 29, 47, -33, -44, -90, 
        -88, -38, 98, 58, 36, 51, -51, -63, -113, 
        -94, -55, -73, 53, -122, -80, -93, 68, -71, 
        -19, 63, 81, -6, 66, 13, 12, 5, 76, 
        -119, -98, -9, 24, 53, 11, -46, 13, 62, 
        26, 82, 30, -84, -54, -65, -82, 51, -61, 
        74, 106, 102, 36, 107, -51, 108, 6, -37, 
        85, -14, -38, 89, -13, 4, -29, -90, -107, 
        23, -15, 11, -43, 80, -88, 62, -19, 16, 
        -67, -16, -89, -35, -71, -17, 1, 13, -31, 
        -77, -96, -93, -55, 60, -79, -97, -44, -84, 
        61, 47, -88, -85, -3, -27, -51, -95, 0, 
        46, 18, 39, 32, 49, 35, -53, -40, -17, 
        -9, -15, -6, 22, 13, 40, -29, -10, 15, 
        -39, -17, -2, -64, -86, -60, -18, -41, -25, 
        9, -18, -12, 18, 1, 34, -5, 2, 3, 
        -4, 22, -2, 5, -14, -23, 6, -17, -1, 
        0, 23, 1, -50, -37, -29, -18, -13, -4, 
        -23, 2, 27, -64, -43, -38, -19, -56, -6, 
        22, -5, -7, 0, 22, 18, 13, -6, 6, 
        4, -17, -27, 37, 20, 16, 30, 67, 37, 
        -3, -35, -19, 23, 27, 16, 3, -25, -18, 
        -12, -11, 3, 4, 23, -13, -13, 4, -16, 
        -18, -43, -50, 36, 38, 21, -42, -13, -35, 
        40, 41, 72, -42, 31, 31, -11, 24, 7, 
        -18, 0, -5, -1, -16, 3, 14, 1, -5, 
        -1, 9, 0, 1, 26, 48, -28, -44, -26, 
        8, 0, -11, 22, 26, 42, -6, -9, 2, 
        7, -21, -41, 39, 21, 34, -33, -19, -14, 
        2, 17, 8, -69, -20, 9, -22, -17, -11, 
        10, 18, -15, 19, 12, -3, -21, 4, -6, 
        -5, -2, 4, -16, 13, -9, -15, -6, -15, 
        12, -5, -14, 22, 49, 33, -44, -47, -18, 
        -38, -1, -14, 29, -19, -52, 16, 33, 27, 
        23, 35, 5, 19, 28, 37, -19, -27, -46, 
        31, 26, 7, -11, 50, 46, -62, -56, -30, 
        33, -1, 10, 1, 25, 8, -10, -27, -18, 
        16, -21, -13, -14, -17, 2, 7, -11, 13, 
        -33, -71, -96, 34, 7, -29, 10, 12, -30, 
        15, 6, 19, 18, -2, 1, 9, 6, 10, 
        -11, -1, 8, -12, 2, 6, -12, 1, 2, 
        -21, 9, 13, 59, -6, -9, 78, 127, 107, 
        19, -14, -39, -46, -36, -36, -34, -61, -47, 
        -23, 5, -41, 19, 51, 36, -9, 36, 0, 
        -33, 10, 23, -36, -30, -42, -13, -26, 1, 
        -49, -52, 8, -4, -25, -20, -50, -26, -28, 
        1, 17, 10, 10, 18, 18, 13, 40, 0, 
        -38, -42, 37, -40, 18, -11, -8, -36, -57, 
        -13, -20, -19, -13, -12, -13, 2, 18, 10, 
        13, 38, 7, 15, 43, 22, 12, 16, 41, 
        24, 9, 18, 24, 1, 40, 21, 31, 6, 
        -8, 16, -7, -11, -14, -12, -7, -5, 5, 
        5, -30, 51, 5, 33, 44, -4, 16, 13, 
        -51, -45, 27, -31, 8, -4, -32, -25, -21, 
        -16, 21, -14, -16, 19, -12, -17, 19, 2, 
        -70, -31, 38, -35, -13, -28, -45, -30, -36, 
        -5, 20, 67, 32, 4, 30, 16, 21, 31, 
        10, 17, 7, 3, 17, -15, 19, 16, 17, 
        -33, -30, 40, -46, -25, -20, -26, -26, -42, 
        -48, -37, 12, -17, -1, -49, -20, -22, 5, 
        -43, -38, 47, -53, -30, -41, -38, -7, -6, 
        -57, -10, 127, -69, 4, -38, 5, -18, -47, 
        -5, 7, 20, -4, -10, -3, 1, -6, 0, 
        5, -8, -8, 2, 17, 1, -9, 12, 14, 
        -50, -53, 37, -26, 7, -41, 17, -18, -47, 
        -8, 28, 45, 6, 5, 19, 34, 12, -2, 
        -49, -19, 19, -58, 20, -27, -29, -20, -1, 
        -48, 6, 42, -44, -11, -71, 5, 5, 23, 
        8, -20, 28, 10, -24, 7, -2, -12, 23, 
        4, -16, -11, 10, 15, 9, -22, -3, 17, 
        5, -91, 25, -15, -19, -8, -28, -32, -33, 
        17, 17, 5, 2, 15, -17, 2, -19, -9, 
        -3, 1, -16, 14, -9, -3, -18, 15, -7, 
        3, -6, 56, 31, 42, 26, 2, 35, 9, 
        -58, -7, 28, -46, 45, 11, -46, -18, -69, 
        -26, -42, 36, -6, -28, -16, -46, -58, -33, 
        -9, 17, -27, 7, -36, -17, 14, 10, 57, 
        6, 35, -37, 9, 23, -40, 10, -2, -29, 
        -6, 45, 38, -34, 41, 25, 37, -24, -18, 
        -7, 44, -16, -14, 25, -47, 28, -28, -33, 
        -21, 26, 9, -25, 23, 22, 20, 8, -14, 
        -4, -69, -33, -30, -67, -15, -20, -59, -41, 
        -9, 6, 26, -40, 29, 14, 14, -23, -59, 
        0, -21, 3, -25, -11, -23, -9, 21, -21, 
        -53, 13, 33, -34, -17, 1, 18, 27, 25, 
        29, 48, -16, 18, -1, -40, 8, -18, 11, 
        -1, 0, 0, -17, -2, 16, -12, 8, 12, 
        22, 40, -49, 46, -10, -60, 21, 9, -1, 
        -28, -52, -44, -101, -41, 10, -37, 54, 60, 
        -8, -11, -3, -7, 6, -20, -9, -12, -3, 
        -9, 55, 8, 29, 34, -54, 0, -37, 11, 
        30, 35, -47, 3, 1, -34, 6, 0, 20, 
        -2, 32, -30, 10, 7, -42, 11, -25, -21, 
        50, 99, 101, 86, 31, 41, 11, -8, 29, 
        14, -17, -24, -16, 10, 1, -14, 5, 12, 
        -16, -14, 9, 20, -22, 10, 6, -6, -4, 
        33, 53, -4, 45, 20, -53, 46, 7, 25, 
        -27, -36, 33, -39, -1, -28, -16, 40, -7, 
        20, 37, -65, -4, 0, -27, -11, 18, 8, 
        -8, 7, -58, 44, 7, -4, -11, -5, 51, 
        -1, -1, -10, -28, -22, -41, -6, -4, -14, 
        21, -23, 10, -3, -24, -7, 4, 19, 25, 
        56, 36, -25, 27, -64, -10, -4, 40, -43, 
        21, -23, -2, -18, 17, -22, -14, -13, -21, 
        -18, -12, -4, -14, -8, 18, -9, 4, -24, 
        -127, -80, 26, -127, -65, -11, -50, 28, 32, 
        14, 108, 78, 82, 79, -45, 35, 7, -49, 
        -5, -15, -40, -20, -56, -78, 19, -7, 25, 
        9, 37, 49, -77, -1, 11, -47, -42, -17, 
        23, 6, 58, -22, 37, 23, -74, -45, -18, 
        -8, -11, -56, -28, -37, -18, -38, 6, 35, 
        -1, -20, 37, -17, 25, 19, -50, -44, -28, 
        28, -19, 21, 19, -2, -10, 2, 18, -16, 
        -12, -30, -32, 31, 4, -22, -4, -25, 37, 
        -17, 2, -65, 15, -38, -60, -41, -4, -8, 
        -29, 6, -13, 2, 6, -29, -3, 31, 9, 
        -24, 22, -18, 12, 24, 30, -36, 28, -8, 
        -32, 31, 50, -9, 0, 80, -85, -50, -43, 
        -18, 5, -7, 12, 0, -25, -5, -12, 20, 
        -25, 19, 16, -21, 25, 83, -92, -50, -35, 
        -40, 34, 33, -22, -17, -48, 25, 31, 79, 
        -10, 16, -25, 24, 8, 7, 13, -21, -13, 
        19, 4, 43, -38, -23, 16, -89, -28, -30, 
        23, 40, 36, 11, 19, 63, -29, -80, -48, 
        15, -7, 28, -26, 28, 57, -25, -40, -42, 
        -35, -12, 38, -127, 70, 36, 109, -42, -70, 
        -1, 17, -20, 19, -26, -5, 16, -21, 5, 
        31, 9, -1, 2, 21, -2, -16, -6, -8, 
        9, 10, 60, -21, 20, 25, -32, -47, -54, 
        -52, -35, -38, 22, 34, 10, -11, -8, 38, 
        -39, 3, 44, -70, -13, -31, -37, -46, -54, 
        -21, 14, 75, -85, 1, 15, -53, -75, -64, 
        11, 29, 48, -6, 4, 53, -82, -64, -61, 
        0, 16, -6, -2, 13, 4, 21, -6, -1, 
        -21, -36, 7, 40, 1, 33, 0, -84, -60, 
        2, 16, 23, 22, 9, 21, -11, 28, -16, 
        -10, 11, 27, -31, 19, -27, 16, 18, 28, 
        -43, -8, -64, -12, -22, 76, 40, 93, 95, 
        -4, 37, -60, -41, -39, 7, -101, -74, -114, 
        33, 39, 11, 1, 42, 91, -44, -42, 41, 
        -19, 39, 39, 2, 23, 3, 30, -45, -36, 
        -11, -25, 21, 6, 2, -2, -11, 4, -39, 
        -18, -36, -3, -22, 5, 7, 25, 44, 26, 
        -44, -22, 10, -6, 19, -4, 15, 20, -13, 
        16, -5, 16, 16, 10, 8, -2, -12, 7, 
        3, 0, -14, 10, -18, 10, -19, -16, -1, 
        -5, -13, -24, 12, 0, 6, 3, 15, 17, 
        -13, -11, 18, -12, 17, 16, -9, -4, -13, 
        -5, -40, 14, -7, 8, 30, 27, 30, -5, 
        -39, 7, 3, -1, 3, -10, 13, -11, -32, 
        1, -5, -9, -18, -12, -18, 6, 11, 8, 
        -63, -33, 5, 8, 14, 2, 10, -21, -36, 
        -8, 33, -9, 3, -25, -7, 8, -20, 4, 
        1, 7, 12, -21, 17, 4, 12, 12, -1, 
        -32, -10, 27, -14, 31, 4, 38, -19, -55, 
        -15, -17, 26, 5, 10, 9, -12, -20, -13, 
        -21, 3, 31, -8, 35, -5, 8, -34, -34, 
        -55, 43, 54, 45, 95, 44, 127, 55, 49, 
        14, 10, -4, -12, -3, 17, 6, -13, 6, 
        -10, 13, -10, 13, -9, -11, 0, 13, -16, 
        -59, -13, 29, -3, 42, 20, 37, 0, -56, 
        -7, -24, -20, -2, -3, -19, -24, 29, 23, 
        6, 21, 1, -3, 26, -5, 19, -29, -33, 
        -15, 10, 15, -3, 24, -15, 23, -29, -50, 
        -34, -17, 16, -7, 3, 9, -18, -6, -19, 
        5, 9, -10, -17, -15, -18, 14, -13, 18, 
        -24, -12, -21, 19, -32, -29, -56, -41, 6, 
        16, -4, 10, 9, 12, -1, 13, 3, -8, 
        -4, 17, -2, 7, -14, 16, -19, -3, -13, 
        20, -1, -1, -14, -5, -14, -27, 41, 22, 
        -77, -59, 0, -32, 41, 71, 84, 46, -12, 
        -52, 1, 6, -30, 14, 14, 0, -22, -37, 
        -99, -79, -97, -58, -8, -104, -117, -105, -70, 
        -60, -64, 40, -11, -108, -108, 99, -45, -116, 
        9, -111, -111, 48, -10, 54, -117, -121, -25, 
        -49, -84, 102, 86, -105, -47, -9, -82, -78, 
        77, -90, 26, -74, 26, 68, 77, 10, -71, 
        45, 23, -118, -38, -62, 63, -79, 84, 19, 
        -98, 90, 110, -56, -51, 2, -117, 86, 111, 
        12, 27, -104, -2, 101, -105, 74, -68, -119, 
        -108, -38, 30, 71, 17, 76, -103, 64, 25, 
        93, -39, -90, -47, 88, -96, 67, -15, -24, 
        -84, 82, -100, 11, -25, -98, 5, -118, -119, 
        -25, -33, 15, 73, -26, -28, 39, -22, -53, 
        -109, 92, -118, 6, 60, 10, 86, -71, -72, 
        5, 82, 61, -94, -112, 30, 42, 103, -24, 
        87, -66, -59, 91, -127, 76, -13, 70, 17, 
        -43, 41, 30, -16, -124, -21, -43, -114, 8, 
        -7, -53, -111, -125, 12, 40, -45, -89, 86, 
        -103, -6, -61, 54, -64, 42, -89, -90, -24, 
        79, 99, 107, -29, 78, 14, -1, -5, 8, 
        39, -28, -121, -24, 70, 6, -92, -111, 105, 
        41, 57, 114, -4, 32, -80, 45, 105, 42, 
        -25, -25, -75, -48, -23, 6, -88, 15, -56, 
        25, -53, -88, 104, 3, 70, 14, -3, 16, 
        -93, 86, 51, 10, 59, 27, 34, 75, -14, 
        24, -77, -66, 8, 57, 95, 54, -86, -10, 
        -7, 110, 45, 32, 0, 86, 62, -26, -79, 
        0, -117, 46, 25, -116, -120, -117, -9, -105, 
        -52, 80, 94, 94, 52, -20, 60, -98, -109, 
        -1, -28, 28, 32, -19, 69, -72, -52, -13, 
        -57, -68, -30, -43, -98, 38, -23, 29, -50, 
        -103, 26, 92, -119, -23, -16, 0, -112, 81, 
        -70, -80, -91, 88, 8, 81, -73, 28, -113, 
        -110, 26, 53, 28, -23, 83, 72, 35, 3, 
        76, 52, -9, 24, -2, -113, -16, 36, 55, 
        -35, -92, -31, 51, -23, -42, -127, 17, -9, 
        -21, 60, 29, -89, 32, -79, -33, 5, -111, 
        56, 68, 73, -1, -49, 73, 90, 12, 47, 
        67, 86, -69, -15, 45, 12, -98, -91, -37, 
        -92, 81, -82, -68, 68, -27, 18, 25, -30, 
        74, -48, -90, 34, -95, -15, 16, -28, 36, 
        -76, -3, -90, 43, 35, -15, 20, -49, -105, 
        -6, 74, 15, 50, 25, 14, 8, -25, 33, 
        32, 71, -38, -19, 95, -45, -58, -31, 1, 
        -119, 16, 83, -41, 61, 65, 55, 73, 76, 
        5, -41, -93, -36, 33, 17, -74, -30, -47, 
        -18, 3, 35, -77, -31, -52, -15, -46, -67, 
        -55, -72, -89, -54, -93, 75, -29, 15, 60, 
        -5, -12, 42, -27, -119, 28, -56, -11, -70, 
        -87, -13, 73, -18, -29, -40, 45, 43, -43, 
        -71, 54, 97, -41, 30, -37, 95, -92, -78, 
        -72, 15, -73, 47, -38, -90, -4, -53, 46, 
        21, 15, -40, -18, -66, -36, -61, 64, -87, 
        20, -4, -65, -22, -97, -61, -5, -4, 24, 
        -39, 35, -78, -84, -121, 47, -77, -99, -9, 
        17, 28, 35, 36, -16, -83, -57, 64, -28, 
        -94, 26, 20, -36, 69, -94, 15, 75, 75, 
        -38, -65, -97, -62, -113, -97, -56, -69, -57, 
        17, -91, -2, -6, 81, -52, 60, -43, -26, 
        -69, 87, -102, -39, 14, 67, 16, -12, 20, 
        -50, -45, 67, -23, -96, 71, -94, -9, 49, 
        14, 63, -65, -39, -87, 26, -41, 24, -64, 
        -82, 82, 32, -127, -44, -83, 36, -8, -92, 
        -95, 46, -103, 70, -115, -98, -25, 66, 70, 
        -110, 75, -50, -2, -94, 14, 4, 49, 39, 
        2, 30, 27, -71, -43, -90, 19, -8, 13, 
        33, 36, 17, -45, 0, -19, -17, -7, 2, 
        -16, 16, 18, -42, 24, 63, -19, -10, -25, 
        2, 18, 42, -20, 7, -19, -10, -30, -27, 
        -19, -12, 5, -16, 18, 3, 15, -13, -10, 
        -13, -21, 34, 10, 13, 15, 20, 25, 22, 
        13, 1, 28, 5, -3, 30, -2, 16, 22, 
        12, -14, 16, 13, 16, -4, -13, 5, -3, 
        19, 14, 42, -11, 29, 24, -18, -17, -7, 
        30, 50, 12, -37, 6, -75, -20, -20, -29, 
        11, 14, -21, -5, 9, -7, 3, 6, 2, 
        27, 47, 42, -19, 9, -72, -4, -47, -22, 
        -35, 13, -38, 9, -6, 50, 6, 38, 23, 
        -2, 15, -16, -23, -4, -4, 5, -3, -23, 
        5, 30, 22, -68, -30, -49, -9, -8, -21, 
        16, 38, -11, -53, -22, -58, -17, -30, -12, 
        30, 39, -1, -22, 5, -44, 3, -23, -8, 
        -97, 14, 84, -58, -11, -33, -5, 37, 7, 
        14, -12, 19, 7, -13, 3, -10, 21, 14, 
        8, -21, 6, 14, 13, -1, 10, -18, 3, 
        -5, 35, 41, -69, -4, -50, 2, -23, 13, 
        44, 12, 6, 26, 0, 1, -10, -21, -18, 
        -25, 7, 17, -70, -34, -72, -17, -9, 23, 
        -1, 18, -5, -79, -53, -69, 22, 6, 33, 
        24, 19, -6, -35, -7, -53, -19, -10, -2, 
        20, -9, -14, 0, -19, 10, -19, 21, -4, 
        19, 24, -83, 65, 13, -127, -72, -75, -20, 
        -20, -5, 2, -8, 3, 20, -19, -2, -14, 
        -13, 8, 20, -19, -12, 3, 3, -20, 4, 
        10, 1, 0, 42, 53, 26, -12, -1, -13, 
        -25, 20, 52, -100, -26, 45, -22, -38, -115, 
        47, 24, 29, -28, -8, -68, -38, -27, -16, 
        -86, -102, -76, -73, 100, -103, -7, -58, -87, 
        66, -51, -107, -71, -70, -73, 97, -32, 47, 
        28, 19, -51, -31, -92, 22, 60, 86, -66, 
        -63, 33, -98, -6, -41, 87, -71, -75, -6, 
        -9, 56, 18, 19, 23, -93, -91, -102, -49, 
        36, -109, -30, -28, 38, 10, 94, -72, -127, 
        5, 24, -73, -2, -107, -95, -1, -110, 51, 
        -99, 14, -28, 83, -92, 62, 26, -46, -104, 
        18, -39, 1, 34, -117, 17, -105, 60, 62, 
        -90, -41, 29, -71, -17, -96, 15, -63, -92, 
        -76, -16, -1, 77, 90, -89, 75, -97, -95, 
        -18, 29, -5, 90, -58, 81, 50, -26, -10, 
        43, 7, -60, -17, 0, 95, -46, 56, -85, 
        -58, -55, -66, 0, 68, 106, -54, -91, -89, 
        29, 40, -81, -61, 34, -66, 32, -117, -6, 
        46, -22, 10, 79, -49, 52, -27, 0, 62, 
        -117, -42, -88, -94, 5, 46, 38, -92, 0, 
        57, 86, -16, -53, 19, 51, 23, 37, -42, 
        -59, 13, 48, 55, -68, -99, -71, 56, -101, 
        71, 37, -87, -100, -21, 58, -22, -90, 89, 
        58, -36, -31, 3, 84, -48, -7, 26, -99, 
        80, -110, -21, 80, 83, -11, -95, 24, 89, 
        67, -86, 72, -107, 95, 56, 16, -20, 93, 
        73, -11, -10, -54, 14, 56, 19, 29, -75, 
        24, 29, -65, -41, 0, -1, -76, -85, -24, 
        22, -108, -49, 85, 58, 54, 48, 84, -80, 
        -67, 95, 87, -29, 96, -48, -17, -62, -28, 
        5, 5, -108, 110, -3, 14, -58, 13, 12, 
        6, -107, 54, 11, 71, -4, 32, -36, -48, 
        82, -91, -106, 90, -93, -95, -83, 86, -57, 
        -10, 17, -7, 36, -105, 99, 79, 44, -54, 
        -31, -71, -110, 95, 68, -22, 18, -2, 73, 
        -11, 18, 38, -21, -23, 9, -67, -24, -31, 
        22, -5, 0, -26, -9, 0, -39, -36, -1, 
        -18, -60, -61, -5, -41, -94, 31, -12, -1, 
        1, 25, -25, 9, 21, -1, -21, -25, -6, 
        10, -8, -4, 0, 14, -13, 6, 9, 3, 
        0, -32, -17, 2, 16, -23, 11, -5, -29, 
        8, -52, -29, -12, -9, -35, 34, -12, -34, 
        6, 7, 17, -10, 10, -4, -1, 17, 13, 
        8, 25, -27, -13, 14, -13, 5, -11, 18, 
        -11, 0, 12, 4, 14, 40, -34, -43, 7, 
        4, -19, -17, -5, -17, -14, -14, -9, 1, 
        -12, 28, -6, -12, 17, 35, -2, -7, -19, 
        20, -4, 91, -2, -1, 17, -16, 13, 5, 
        -9, 19, -18, 8, -15, -8, 1, 20, 1, 
        5, 24, -6, -27, -22, 11, -33, -23, 7, 
        5, 9, 14, -32, 3, 6, -8, -36, 21, 
        12, 15, -23, 8, 16, 14, -5, -38, -5, 
        33, -34, -75, 22, -52, -127, 20, 94, -5, 
        22, 10, -4, -7, -2, 17, -10, 12, -20, 
        0, 11, 3, -11, -15, 19, 10, 4, 12, 
        18, -4, -9, -20, -36, 7, -30, -12, -4, 
        7, 26, -3, -31, -11, 10, -1, -12, 29, 
        -17, 42, 35, -41, -35, 17, -20, -22, -19, 
        0, 29, 9, -19, -35, 7, -20, -11, -5, 
        3, 23, 16, 9, -5, 13, -30, -43, -20, 
        -7, 3, -8, -5, -17, -17, -4, 18, -15, 
        37, 42, 25, -25, 6, 99, -17, -14, 34, 
        7, -8, -1, 14, -1, -21, 16, -1, 7, 
        -7, 9, 17, -5, 5, -12, -8, -16, 8, 
        61, 57, 21, -12, 23, 27, -13, -13, 30, 
        -26, -50, -3, 6, -37, -58, -22, -32, -10, 
        32, 47, -7, 8, 11, 27, -21, -41, 54, 
        -15, -6, 1, -32, 10, 1, 15, 6, 0, 
        -8, 18, 17, -38, 0, -9, -28, -5, 0, 
        27, -23, 45, 30, 30, 13, 30, 68, 49, 
        14, 7, -19, -30, 8, 40, -49, 18, 25, 
        -6, -31, 10, -5, 15, 4, 11, -25, 18, 
        19, -28, -25, 28, -2, 25, 12, -22, -18, 
        -15, -7, -36, -8, 3, 57, 1, 28, 20, 
        30, 9, -8, 28, 8, 18, 15, -29, 20, 
        31, -51, 23, -42, -15, 5, -65, -15, -29, 
        -20, 2, -7, 0, 0, 11, -16, 63, 13, 
        -1, -19, -16, 8, -2, -4, -9, -29, 8, 
        15, 60, 5, -87, 40, 11, -11, 22, -13, 
        -20, -32, -10, 15, -101, -71, 8, -69, -104, 
        -25, 28, -21, 26, 1, 1, 4, -32, -1, 
        -49, 5, 36, -60, 12, 28, 2, 56, 25, 
        -5, 24, -1, -52, 4, 1, 6, 39, 52, 
        -4, 15, 0, -44, 2, 34, -17, 39, -15, 
        34, -5, -41, -19, -6, 8, 105, 75, -12, 
        5, 33, -17, -18, 32, 33, -35, 24, -4, 
        -3, -20, 13, 26, 33, -14, 0, -27, 17, 
        -62, -33, 0, -48, 42, 37, -9, 26, 11, 
        4, 20, -23, 84, -30, -50, 13, -50, -18, 
        27, 11, -3, -99, 38, 21, -31, -5, 36, 
        -32, 42, 31, -62, -4, -37, 42, 56, -31, 
        -24, 14, -3, 4, 6, 24, 6, 30, 8, 
        0, 26, 5, -22, -34, -31, -7, -15, -27, 
        78, 121, 61, 57, 85, 42, -2, 48, 71, 
        0, -32, -6, 9, -2, 18, 14, -33, -16, 
        34, 2, 7, -3, -24, 15, -31, 26, -23, 
        13, -71, -82, 49, -92, -127, -19, -101, -92, 
        -43, -21, 82, -47, 52, 56, 22, 104, 49, 
        24, 54, -10, 45, 26, 14, 39, -6, 5, 
        -28, -98, 86, -62, 81, 97, 69, 57, -74, 
        -39, 14, -53, 58, -103, -99, 27, -20, 86, 
        68, -19, -85, -24, 84, 68, 81, -109, -108, 
        -18, -74, 63, 76, 87, -106, 34, -73, -110, 
        75, 7, -101, -95, 99, 77, -87, 51, -85, 
        -2, 21, -61, 41, -108, 44, 66, -94, 27, 
        -88, -104, -42, 55, -34, -43, 3, -48, 85, 
        83, -40, -18, 64, -30, 84, 97, 102, 41, 
        -62, 3, 5, 27, 50, -20, 29, 11, -88, 
        -55, -48, -11, 81, 11, 41, 55, -23, 107, 
        -7, 48, -110, 63, -60, -88, 56, -6, 55, 
        -2, -73, -106, 3, -101, -27, 42, 47, -41, 
        -87, 0, -96, -18, -13, 44, -39, -96, 90, 
        34, 90, 3, 61, -3, -99, -84, -89, 62, 
        0, 18, -105, 88, -14, 52, -83, 61, -102, 
        -92, 18, 18, -72, 43, 50, 62, -73, -29, 
        88, -41, 52, -115, 12, 37, -120, -16, 86, 
        9, -40, -95, -2, 101, -60, 68, -11, 96, 
        24, 9, -69, -111, -8, -5, 91, -33, -76, 
        81, 9, 16, -22, -89, -90, -107, 3, -83, 
        62, 53, 61, 4, -58, -29, -95, 88, -89, 
        3, 22, -44, 59, -37, -110, 66, 52, -29, 
        -37, -21, -30, -127, -52, 103, 83, -49, -26, 
        35, -45, 56, 45, -86, 121, -17, -80, 87, 
        -104, -10, -12, 80, 62, -17, -41, 33, -86, 
        -53, 9, 0, 1, -86, -38, 29, 63, -88, 
        -76, -1, -22, -104, 88, -106, 102, -93, -83, 
        19, -107, -108, 94, -70, 13, 55, 85, -76, 
        -48, 27, -39, -35, 103, 101, -77, 64, -5, 
        -111, 27, 22, -30, -18, 47, -86, 19, 4, 
        29, -44, 68, -78, -33, -94, -46, 109, 99, 
        -27, -11, -93, -14, 20, -118, -89, -51, -39, 
        -59, -30, -76, 79, -9, -60, 55, -49, 8, 
        -91, 41, -47, 37, 20, -50, 31, 52, -98, 
        19, 9, -36, -127, -4, 34, -95, -37, -59, 
        -76, 61, 46, -92, 22, 61, 5, -76, -77, 
        23, -28, 12, 80, -61, -11, 17, -38, -41, 
        -42, -10, 53, 35, -59, -99, 20, -83, -27, 
        -84, 3, -21, 53, -36, -75, -89, 16, 51, 
        89, 87, -73, -85, 85, 13, 12, 85, 64, 
        -81, -32, -99, -22, 21, -30, -84, 7, -63, 
        -92, 32, -104, 21, -74, 18, -62, 8, 27, 
        84, 9, -76, -2, 45, 34, -74, -34, 85, 
        -51, 82, -59, -93, 9, -3, 18, 34, -67, 
        1, -46, -93, -119, -78, -97, 29, -4, 16, 
        17, -32, 18, 2, 39, -83, -22, 3, -68, 
        14, 70, 4, -3, 38, -26, 23, -27, -9, 
        -77, 61, 74, -69, -6, -65, -27, -121, -115, 
        51, 63, -75, -65, 59, -88, -91, -51, 17, 
        -14, 69, 91, 37, 89, 59, 0, -66, -74, 
        86, -29, 28, 62, 77, 43, 80, -13, 63, 
        -41, 9, 58, 27, -93, -66, -7, -7, 54, 
        -47, -80, 64, -29, -98, -37, -67, -95, 26, 
        -58, -38, 40, 51, -28, 60, 3, -80, 5, 
        81, 18, 2, -4, 57, 33, -8, 20, -37, 
        44, 55, -60, 59, -33, -41, -4, 51, -88, 
        -94, 16, -46, 34, -96, -89, -4, -119, 48, 
        -70, -40, 38, 46, 15, 4, -64, 66, 92, 
        10, -9, 9, 39, -80, -46, -1, -12, 13, 
        93, 28, -5, -85, -16, 1, 85, -86, 1, 
        -83, -88, -90, 45, -11, -51, -39, -26, -21, 
        27, 8, -64, -15, -106, 27, 41, -91, 48, 
        -11, -84, -71, -8, 14, 73, 49, -68, 66, 
        84, -104, -19, 71, 14, -74, -83, -35, 2, 
        -75, -25, 33, 67, -4, 82, -36, 50, 55, 
        3, -60, -19, -82, 52, -97, -41, -40, 4, 
        -100, 69, -30, -102, -102, 71, -102, -11, 78, 
        -28, -124, -46, -75, 87, -90, -1, -47, 14, 
        34, 12, -18, -64, -37, 79, -94, -26, -82, 
        15, 59, 63, -52, -112, 11, 61, -68, 87, 
        -67, -10, -72, -11, 10, -123, 64, -10, 31, 
        -71, -35, 64, 17, -34, -26, 8, -82, -100, 
        -103, -90, 5, -72, -24, -60, -17, 82, -39, 
        11, 80, -58, 20, -106, 42, 103, -90, -118, 
        -18, -9, 6, -44, -111, -100, 61, 73, 9, 
        -27, 54, 78, -23, -7, 63, -5, -32, 44, 
        -55, -19, 54, -75, 76, 10, 31, -58, 55, 
        36, 111, -83, -74, -79, 38, -73, -16, 45, 
        -51, -28, -20, -61, 52, 21, 22, 77, -35, 
        70, 86, 69, -78, -111, -58, -7, -100, -99, 
        64, -54, 37, -16, -15, 90, -113, 8, 12, 
        44, -85, -40, 55, -58, 40, 43, -113, -101, 
        -1, 79, 29, -63, 32, -99, 33, -50, 48, 
        -21, 96, 35, 56, -65, -88, -21, 11, 44, 
        -2, -92, 48, -80, -48, -91, -58, -105, -117, 
        -55, 80, 38, 80, -31, -74, -100, -56, -72, 
        -114, 4, 73, 15, -75, -36, -61, 58, -101, 
        -17, -99, 50, -2, -115, -102, -1, 63, -22, 
        -124, 52, -44, 34, 49, -34, 10, 88, -48, 
        -58, -6, 89, -58, 84, -23, 83, 107, 93, 
        -112, -125, -85, -71, 100, -79, -40, -6, -15, 
        45, 88, -6, 32, 49, 22, -106, -26, -21, 
        25, -107, -61, 99, 107, 93, 4, 64, -106, 
        -90, 28, 70, -10, -127, -117, -65, 87, -111, 
        -17, -2, -81, 100, -110, -68, -79, 61, 33, 
        -79, 63, -2, 33, 81, 37, 75, -50, 35, 
        -89, 54, -39, -21, 9, 6, -72, 29, -91, 
        -25, -3, 57, 20, 39, -100, -44, -52, -73, 
        12, -55, 59, 38, 51, -53, -37, -106, 36, 
        -78, -60, 45, 58, 10, 74, -89, -67, 48, 
        53, 70, 87, -58, -51, 32, -7, -70, 76, 
        -87, -44, -112, -94, 77, -90, 67, 12, -14, 
        -4, 16, -75, -100, -26, -20, -8, -67, 90, 
        5, 49, -85, 54, 95, 19, -100, -90, 58, 
        67, -74, -32, 67, -40, 79, -93, 54, -22, 
        36, -47, 40, 2, 63, -69, -105, 46, 80, 
        -23, 33, 27, -42, -30, -9, 36, 0, -97, 
        19, 56, -115, -124, -57, -127, -91, -58, 67, 
        -23, 4, -2, 90, -45, 51, -96, -106, 27, 
        87, -35, -57, 98, 33, 91, -42, 93, 74, 
        65, -114, 3, -91, -71, 40, 77, 66, -3, 
        82, -18, -27, 76, 80, 51, -93, -76, -80, 
        72, -30, -109, 46, 27, -48, -11, 16, -92, 
        78, 76, 24, 65, -2, -22, 99, 85, -93, 
        90, -83, 105, -1, -42, 58, -14, 93, 75, 
        -89, -106, 95, -72, -6, -37, -77, 19, 107, 
        -59, 29, 22, 17, -55, 60, -89, 23, 16, 
        58, -108, -9, -77, 92, 61, 53, -95, 44, 
        -116, 3, -10, 3, -8, -111, -4, 44, -19, 
        -10, 78, -29, -105, 94, -82, 7, -89, 72, 
        -35, -15, -14, 45, -64, 14, -88, 86, 86, 
        2, 49, 80, -12, -97, 44, 16, -58, 99, 
        -8, 82, -26, -46, 63, -74, 57, 94, -43, 
        -91, -98, 98, 107, 37, -52, -44, -80, -28, 
        -74, 3, 53, 17, -6, -51, -94, 45, -96, 
        -81, 86, 69, -104, 42, 37, -41, 86, -56, 
        73, -32, 28, 0, -88, -52, -43, -60, -116, 
        75, 58, -104, -51, 48, 5, -72, -58, 86, 
        1, 23, 12, 15, 14, -5, 46, 5, 50, 
        1, -26, -14, 10, 42, 5, 10, -11, 53, 
        -29, -42, -25, -87, -63, -95, -51, -47, -82, 
        -14, -29, 27, 0, 8, -3, 29, 49, 31, 
        0, -13, 6, 5, -4, 32, 18, -5, 19, 
        43, 5, -16, 19, -14, -20, -25, -53, -53, 
        22, -36, -15, -57, -91, -85, -85, -96, -43, 
        9, -15, 8, -4, -3, -16, -32, -4, -33, 
        -29, -31, -59, 5, -8, 46, 31, -22, 42, 
        -11, -43, -32, 38, -16, 0, 19, 48, 1, 
        14, -1, -28, 6, -27, -2, 17, 21, 27, 
        -57, -9, -4, 23, 15, 27, 54, 5, 2, 
        88, 75, 21, -12, -70, -89, -19, 16, -59, 
        -22, 5, 0, -4, -9, 31, 8, 14, -6, 
        20, -20, -6, 51, 46, 43, 72, 3, 3, 
        18, 19, 10, 32, 33, -6, 58, 39, 18, 
        -39, -31, 1, -6, 21, 15, 25, -10, 55, 
        26, 62, 38, 68, 41, -16, -18, -34, -65, 
        14, -34, 2, 26, 13, -29, -4, 29, -11, 
        29, -6, 14, 18, 4, 13, 28, 1, 23, 
        -26, -7, 13, 6, 21, 49, 24, 57, 19, 
        10, -51, -26, -64, -98, -55, -94, 0, -20, 
        25, 11, 50, 29, -23, 25, 6, -2, -1, 
        39, 61, 17, 15, 31, 14, 84, -16, 21, 
        -39, 31, -21, -10, 52, 36, 58, 16, 42, 
        15, -31, 2, 0, -26, 24, 22, 17, -33, 
        -16, -12, -71, -44, -36, -2, -86, -108, -24, 
        34, -34, -23, -19, 12, -4, -27, 24, 22, 
        15, 28, 4, -8, -5, -15, 22, -10, -1, 
        32, 22, -94, -127, -108, -72, -86, -37, 45, 
        -29, -34, -58, -14, -44, -45, -18, -31, -26, 
        -27, -28, -24, -51, 1, 54, 5, 10, 5, 
        24, 12, -28, -25, -16, 10, -1, -11, 27, 
        -2, 26, -41, 0, 30, 11, -10, 17, 7, 
        -25, -35, 20, -24, -82, -40, 7, -19, -17, 
        -11, -11, -32, -12, 16, -36, -36, 6, 13, 
        -12, -11, -3, 15, -13, -17, 14, 0, -4, 
        -19, -63, -21, 8, -77, -33, 23, -6, -47, 
        -41, -50, 2, -12, -65, -27, -21, -37, -57, 
        -19, 16, 13, 14, 15, 10, 11, -5, -15, 
        11, -13, -49, -24, 10, -28, -14, 16, 17, 
        3, 35, -56, -17, 32, 8, -6, 21, 15, 
        7, -13, -13, 18, 7, 1, -2, 2, -2, 
        30, 32, -27, -6, 48, -5, -4, 7, 3, 
        -31, -9, 31, -63, -38, 33, 2, -21, -36, 
        1, -18, -14, -17, 6, -3, 9, -15, -1, 
        8, -1, -10, -26, -4, -16, 0, 19, -7, 
        30, 30, -46, -23, 32, 0, 7, -5, 5, 
        25, 13, -20, -4, -11, -4, 11, 18, 18, 
        -27, -13, 44, -29, -62, -51, 39, -7, -47, 
        -13, 18, -12, -1, -3, 15, 16, 4, 9, 
        -16, -17, 15, -17, 7, 4, 4, 4, 11, 
        26, 22, -22, -2, 17, 7, -17, -4, 20, 
        15, -11, -22, 12, -9, -34, -11, 3, -2, 
        17, 31, -5, -38, 35, 48, -3, -17, 14, 
        -2, 14, -30, -10, 4, 8, 20, -15, 6, 
        20, -4, -10, -9, 2, 13, -16, -13, -5, 
        -4, -18, 11, 18, 12, -1, -9, 13, 8, 
        75, 108, -39, 40, 127, 36, -35, -8, 4, 
        13, 10, -1, 18, 10, -18, 13, -14, 14, 
        4, -3, 17, 5, -11, -9, 2, 6, 4, 
        -6, -66, -41, 15, 13, -18, 12, 5, 19, 
        -8, 33, 43, -80, -37, -2, -45, -45, -36, 
        35, 28, -67, 17, 32, -1, -5, 4, 31, 
        0, 25, 36, 33, -21, -35, 7, 4, 23, 
        9, 8, 7, 29, 6, 27, -14, -28, -39, 
        -12, 7, -65, -37, 8, -56, -17, 9, -13, 
        -12, -21, 9, 47, 36, 3, 9, -5, 11, 
        27, -24, 6, 4, -22, 1, -17, 15, 2, 
        -46, -40, -27, -50, -37, -12, -8, -9, 17, 
        -18, -27, -49, -3, -19, -10, -1, -5, 17, 
        21, -26, -18, -11, 12, 20, 9, -18, 4, 
        22, 26, 18, 37, 56, 50, 18, -6, -22, 
        -1, -7, -1, 20, 13, -6, -17, -54, -45, 
        -2, -6, 26, -27, -9, 6, 6, -11, -13, 
        17, 24, 5, 3, 0, 18, -46, -23, -10, 
        70, 43, 99, 16, -18, -17, 44, 116, 38, 
        -2, -11, 19, -16, -17, -23, 22, -21, -6, 
        -19, 12, 8, 20, 16, -5, -19, -55, -6, 
        -6, 5, 21, 21, 36, -4, -43, -52, -32, 
        -2, 10, 26, 19, 24, 2, -1, -31, -16, 
        12, 28, 14, 105, 57, -57, 53, 88, 127, 
        -10, 25, 17, 10, 21, 8, 20, 22, -10, 
        -23, 1, 6, -15, -10, -26, 21, 21, -9, 
        -8, -3, 24, 1, 25, -39, -39, -53, -23, 
        -2, 21, -33, 2, 43, 48, 32, -20, -16, 
        14, 54, 7, -10, -46, 6, -18, 18, -3, 
        -18, 28, 48, 22, -37, -47, -8, -36, 15, 
        16, 20, 19, -4, 8, -13, -14, -44, -29, 
        25, -13, -14, 11, 8, 19, -15, -19, -18, 
        58, 4, -31, -45, 7, 23, 32, -27, -37, 
        0, 17, 11, 28, 12, 8, -9, 20, 13, 
        -2, 20, 4, -6, 16, -5, -23, -26, -17, 
        24, -8, -27, 29, 81, 72, 63, 29, 27, 
        4, -36, -27, 26, -5, -35, -2, -32, -24, 
        7, 20, 30, 19, 36, 38, -21, -21, 1, 
        -43, -62, -35, -83, 25, 62, 81, 75, 9, 
        -27, -12, 22, -15, -20, 33, -22, 36, 28, 
        24, -12, 3, -7, -15, -90, -61, -45, -12, 
        -2, -1, -19, -61, 1, 23, 13, 18, 53, 
        22, 15, 12, 0, 27, -1, -4, 8, -13, 
        -14, -29, 27, -2, -10, -26, 12, -19, 12, 
        20, -2, 39, 12, -40, -21, -36, -55, -33, 
        11, 2, 1, -10, 6, 10, 6, 20, 11, 
        23, 20, 20, -26, -35, 16, -20, 63, 45, 
        -24, -17, 4, -8, -19, 45, 1, 19, 13, 
        16, 11, 24, -5, -11, 26, 26, 25, 20, 
        1, -13, -5, -43, -29, 49, -21, 1, 18, 
        -7, 18, 31, -22, 25, 21, 79, 57, 4, 
        0, -23, 24, 23, -22, -8, -19, -30, 17, 
        -41, -13, -47, -63, -16, 31, 9, 56, 20, 
        0, -6, 18, -33, -5, 9, 25, 28, 25, 
        -37, -36, -8, -62, 13, 24, 22, 15, 47, 
        -34, 17, -100, -103, -43, 45, 107, 120, 127, 
        -29, 6, 7, 22, -11, 4, -11, 12, -4, 
        22, -17, -19, -17, 29, 15, 10, 7, 29, 
        -53, -48, -60, -71, -3, 57, 15, 20, 51, 
        22, 27, 2, 7, -45, -29, 16, 31, 26, 
        -6, -23, -35, -36, 9, 29, 55, 14, -22, 
        -32, -46, -29, -55, 40, 38, 66, 64, 9, 
        -16, -44, 0, -12, 15, 21, -17, 13, -21, 
        4, 21, -5, 10, 22, -14, -18, 0, -20, 
        18, 4, 27, 5, -43, -81, -38, -47, -71, 
        2, 15, 18, 17, 18, 1, 5, -16, 18, 
        -27, 26, -23, 19, -2, -7, -26, 23, -9, 
        28, 54, 32, 15, -5, -82, -27, 58, 24, 
        -65, -13, -65, -110, -126, -86, -64, 44, -33, 
        -8, 32, -23, -11, -16, 32, -24, 47, 21, 
        33, -4, -74, 52, 11, -65, 8, -67, -69, 
        22, 6, -16, 28, -20, -8, 15, -30, -3, 
        -16, -1, 39, 13, 64, 17, 32, 60, -8, 
        23, -23, -19, 0, 51, -38, 40, 24, 19, 
        6, -10, 32, 18, -4, -11, 18, 0, 9, 
        12, 42, 2, 42, 20, 37, 7, 35, 36, 
        11, 25, -15, 37, -4, 40, 46, 5, 3, 
        -19, 4, 7, 12, 26, -26, -10, 0, 0, 
        -10, -8, -28, -51, -41, -52, 17, 4, -29, 
        8, -29, -24, 78, 13, -9, 96, -24, -46, 
        2, -21, 9, 25, 21, -1, 9, -15, 29, 
        16, -39, -71, 50, -30, -11, 63, 34, -28, 
        -31, 9, -45, -105, -25, -38, -76, -84, -32, 
        -12, -29, -10, -1, 9, -15, -27, 28, 26, 
        35, 28, -61, 60, 20, -66, 85, -13, -40, 
        40, 5, -55, 101, 30, -63, 63, -27, -19, 
        61, -6, -19, 55, -24, -58, 76, 6, -38, 
        -64, -126, -70, -27, -79, -76, 10, -102, 26, 
        9, 0, -11, 23, 13, -19, -27, -26, 1, 
        11, 26, -26, 0, -3, -12, -18, -26, 14, 
        45, -29, -68, 39, -41, -25, 106, -23, 11, 
        -34, 16, -24, -53, -21, 3, -15, -56, -1, 
        8, -33, -25, 80, 25, -75, 46, 37, -35, 
        25, -37, -42, 26, -50, -99, 26, -41, 1, 
        38, -2, -9, 59, -8, 1, 32, 30, -34, 
        1, -30, 1, -17, 1, -26, 6, 26, 1, 
        57, 18, -11, 95, 95, 58, 53, -98, 100, 
        -21, 20, 21, 33, 25, -8, 14, -9, 22, 
        -6, -1, -33, 10, 7, -9, -7, -22, -29, 
        -58, -42, -6, -127, -48, -49, -93, -100, -23, 
        -11, 42, -7, 60, 87, 2, 31, 104, -34, 
        -27, 3, -73, 28, -10, -39, -5, -57, -1, 
        -109, -58, -45, 3, -11, -6, 81, -112, 72, 
        -23, 61, 79, -77, -118, -50, -28, 116, 37, 
        -77, -66, 74, -124, 121, -102, 61, 65, 30, 
        71, 100, -57, -4, 106, -3, -8, -12, 20, 
        -112, 119, 104, 102, -67, 78, 21, -112, -95, 
        62, -98, 125, 125, 36, 22, 99, -11, 95, 
        40, 3, -3, -80, 24, -56, -7, -109, -54, 
        -110, -6, 7, -47, -61, -18, 15, 105, -84, 
        -12, 29, -115, -56, 19, 63, -26, 81, -29, 
        32, -58, 7, -111, -31, 26, 76, -24, -109, 
        102, -89, -96, -6, -108, -72, 85, 17, -100, 
        16, -90, -25, 120, -90, 27, -25, -38, 74, 
        -100, 6, 38, -7, -90, -123, -99, -79, -87, 
        70, 53, -20, -78, -45, -15, -38, -1, -111, 
        27, -22, -84, 66, 108, -77, -118, -127, -122, 
        41, -44, -125, 13, 125, -5, -49, -6, -6, 
        37, -49, 28, -101, -4, 19, -73, 86, -109, 
        -120, 107, 115, -50, 15, -39, -103, -123, -47, 
        126, 12, -14, -46, 73, 22, -36, 84, -3, 
        -84, 122, 27, 2, 118, 32, 4, 18, -99, 
        -125, 127, 122, -41, 118, 31, 41, -62, -105, 
        -72, 12, 15, 91, 100, -55, 83, -78, 11, 
        -104, 57, 2, -81, -21, -14, -33, -56, 31, 
        99, -53, -7, -121, 59, 36, -46, -29, -85, 
        -105, -35, -112, 50, 40, -3, 35, 68, -6, 
        44, -97, -37, 10, 111, 111, -12, 96, -9, 
        -16, 9, -19, 22, 102, 33, 118, -75, 50, 
        -107, -48, -13, 11, -88, -58, 42, -7, -99, 
        105, 121, -90, 51, -39, 55, -53, -43, 50, 
        -111, -6, 49, 106, -92, 66, 6, -12, 110, 
        67, -15, -122, 105, 37, -116, -49, 109, 37, 
        -91, 67, -18, -61, -4, 110, 100, -122, -66, 
        -2, 40, -12, -28, -58, -34, -59, 55, 86, 
        22, 52, 18, 30, 5, -58, -57, -29, -7, 
        -14, -25, -35, 4, 43, 14, -21, -11, -28, 
        -23, 54, 40, 39, 33, -45, -43, -61, 2, 
        24, 20, -20, 9, 10, -24, 20, 17, 5, 
        -40, -48, -29, -2, -6, 30, 39, 8, 15, 
        -8, -44, -10, -32, 29, 36, -15, 38, -19, 
        -20, 27, 12, 27, 26, -4, -1, -13, 7, 
        6, 42, 71, 59, 66, 1, -31, -35, 1, 
        31, 27, 11, 3, 6, -54, -62, -11, 3, 
        -25, -15, 28, -23, -28, -21, -24, -22, -17, 
        23, 11, 59, -23, -38, -45, -67, -1, 0, 
        -40, -18, -54, 21, 7, 25, 62, 50, 59, 
        -3, -12, -42, 3, -9, -13, -11, 0, -8, 
        31, 17, 53, -12, -39, -64, -29, -22, 35, 
        1, 3, 42, -15, -34, -24, -64, -13, 43, 
        -4, 55, 65, 6, -23, -66, -72, -19, 23, 
        -10, 69, 50, 34, 16, 60, 9, 87, 113, 
        27, 11, 19, 19, -23, 25, -8, -29, -11, 
        -7, 21, -29, -20, -6, 18, 21, -11, 11, 
        2, 25, 58, 11, -25, -27, -73, 3, 14, 
        -23, -40, 8, 19, 42, -19, 15, -14, -24, 
        9, 23, -4, -5, -58, -63, -58, -12, 56, 
        16, 21, 30, -36, -69, -49, -24, 47, 39, 
        17, 7, 17, 22, -39, -46, -56, -25, 29, 
        20, 16, 19, 27, 19, -23, 4, -16, 28, 
        -16, 15, -30, -2, -67, -120, -75, -75, -92, 
        8, -13, -27, 18, 8, 20, -2, -15, 3, 
        -28, 12, -21, 29, 26, -1, 1, 8, 1, 
        -90, -14, 30, 70, 91, 69, 15, -14, -2, 
        6, 24, 72, 7, 20, -70, -72, -127, -124, 
        -5, 2, 59, 15, -5, -52, -114, -82, 20, 
        -77, -95, 102, -38, -37, -120, -104, -7, -125, 
        80, 41, 3, -57, 94, 81, -36, 61, 106, 
        -83, 78, -55, 4, -76, -79, -22, -107, 68, 
        109, -83, 36, -73, 7, 95, 68, 65, 10, 
        15, -53, -16, 112, -52, -96, 74, -37, 42, 
        13, -8, -26, -114, -55, 79, -105, 85, -101, 
        -121, 53, 72, 27, -1, -97, -7, 54, 48, 
        -57, 105, -43, -12, -27, -119, -76, -100, 103, 
        -118, -91, -117, 54, 78, -79, -114, -65, -81, 
        4, 18, -20, 85, -58, 61, 45, -44, -43, 
        -54, 79, 4, -31, 58, 14, 104, 25, 46, 
        95, -50, -89, 40, 75, 35, -6, -127, -68, 
        72, -109, -111, -42, 18, -84, -102, -5, -92, 
        -9, 70, 88, -111, 116, 93, -79, -85, 27, 
        -40, -100, -95, -67, 54, -23, -43, -41, -77, 
        21, -87, -52, -75, 11, -11, -17, -37, -127, 
        -121, 111, -88, -20, 57, -9, -25, 94, 47, 
        -14, 78, 72, -8, 76, 39, -81, 7, -21, 
        -57, 90, 82, -94, 58, -119, -66, 25, -61, 
        -97, 96, -61, -103, -4, 10, 54, 13, -28, 
        69, 8, 96, -33, 100, 60, 24, 77, 59, 
        57, -11, -83, 59, 47, -117, -6, -123, 103, 
        -6, -9, -22, 6, -115, -24, 108, -7, 105, 
        -78, -90, -16, -11, -61, -8, 65, 82, 17, 
        45, -46, -81, 9, 14, 107, 43, -78, -109, 
        -109, 80, 110, 3, 18, -94, 35, -67, 107, 
        35, -49, -74, 47, 33, 68, 20, 79, -117, 
        -107, -87, 42, -77, -109, -73, -33, -111, -115, 
        116, -10, -41, 44, -40, 27, 7, 91, -99, 
        90, -9, -15, -32, 78, 112, -99, -57, -39, 
        61, -36, -73, 39, -42, -32, -48, 38, -120, 
        -109, 25, 38, -113, -65, 42, 96, 6, -18, 
        -11, 38, 48, 26, 18, -33, 21, 15, -37, 
        -38, 1, 36, 11, 11, -7, 28, -7, -12, 
        -92, -91, -9, -47, 24, 46, -16, -42, -4, 
        -12, 5, 38, 34, 34, 12, 15, 16, -18, 
        -26, -10, -18, -8, -18, -24, 0, 2, -7, 
        -40, -29, -88, -28, -52, -6, -90, -122, -85, 
        -72, -64, -69, -16, 16, 22, -38, -28, -37, 
        11, 21, -24, 6, -4, 22, -25, 3, -23, 
        -36, -15, 60, -20, 30, 0, -11, -29, 4, 
        -3, 25, 5, 23, 11, -11, 24, -13, -27, 
        22, -18, 17, -2, -20, -13, 3, -20, 17, 
        -62, 4, 17, 24, 7, -28, -6, 2, -19, 
        74, 69, -59, -43, -103, 37, -105, 5, -27, 
        10, 3, 6, -3, -20, -16, -30, 14, 23, 
        -6, 32, 24, 23, 24, -45, 38, -3, -29, 
        -22, 8, 26, 35, -7, -40, -6, -35, -31, 
        -40, 17, 40, 18, 25, -29, 21, -36, -4, 
        8, 72, 71, 106, 127, 73, 40, -6, 42, 
        -16, -24, 28, -7, 22, 3, 11, 5, -17, 
        15, 8, -26, 5, -16, 5, -17, -4, -27, 
        -23, 42, 31, 35, 25, -2, 23, -5, -1, 
        -39, -4, -8, -65, -18, 13, -21, -5, -22, 
        -9, 32, 8, 8, 9, -41, -2, -3, -13, 
        5, 62, 47, 19, 17, -38, 42, -23, -11, 
        -35, -3, -19, 9, -15, -32, -7, 23, -59, 
        7, 4, -17, -18, -12, 20, -6, -21, -24, 
        -58, -6, 24, -32, -78, -70, -23, -5, -33, 
        -19, 12, -14, -7, 15, -27, -12, 22, 3, 
        -15, 20, 20, -11, -12, 14, -22, -23, -27, 
        -10, -53, -17, -79, -42, 17, -96, -44, 1, 
        -76, 14, 81, 61, 125, 39, 66, 33, 61, 
        -29, -7, 72, -15, 30, -49, 38, -24, -19, 
        44, -1, -24, 22, 42, 22, 2, 22, 48, 
        15, -52, -40, -9, 17, -10, 5, 1, 7, 
        -4, -21, -18, -15, -52, -11, -47, -69, -41, 
        -25, -14, -45, -13, -12, 10, 17, 32, -15, 
        -10, -12, 24, 10, -21, 9, 11, 24, -19, 
        -31, 5, -9, -37, -38, 4, -62, -75, -34, 
        7, -3, -9, -28, -54, -14, -32, -61, -38, 
        -25, -1, -11, -13, 5, 25, -15, -26, -3, 
        5, -34, 19, 29, -11, -1, 33, 48, 1, 
        -2, -68, -63, -6, 19, -40, 34, 19, 19, 
        -9, 19, -27, 12, -10, -26, -11, 15, -10, 
        -9, -35, -60, 37, -12, -27, 12, 24, -11, 
        16, 24, 19, 30, 31, 52, -13, 1, 18, 
        2, 26, 11, 6, 28, -15, -2, -7, 18, 
        -2, -17, -65, 35, -22, 14, -10, 27, 33, 
        -13, -16, -69, 16, 30, 0, 29, 40, 17, 
        -11, -10, -63, 13, 0, -17, 10, -9, 16, 
        7, 53, 57, -36, -70, -21, 39, -55, 2, 
        13, 9, 2, -22, 20, -11, 26, -25, 13, 
        -15, 13, 23, 26, -23, -24, 6, -16, 24, 
        -24, -24, -64, -8, 11, -36, 25, -18, 16, 
        4, -33, 40, 27, 7, -33, 48, 21, 8, 
        30, 10, -57, 17, 16, 27, -5, 24, 60, 
        22, -14, -51, 11, 21, 20, -12, 12, 44, 
        13, 4, -55, 38, 29, -15, 9, 13, 13, 
        26, 9, -22, 14, -27, 16, 19, -8, -6, 
        20, -41, -38, 53, 65, -73, 40, 127, 16, 
        10, -3, -14, 7, 12, -19, -29, -10, 9, 
        12, 18, 18, 3, 11, -25, -16, 19, -15, 
        -16, -2, 26, 22, -29, 14, 30, 58, 8, 
        46, 25, -16, -18, -62, 26, -2, -30, 29, 
        30, -54, -36, 58, 2, -61, 46, 55, 36, 
        -88, 77, -20, -29, 1, -21, -14, -37, 45, 
        75, -15, 84, 31, -69, -45, -111, 54, -100, 
        -65, 20, -65, 14, -8, 40, -23, 5, 77, 
        76, 90, 83, -81, 93, -88, 60, 47, -98, 
        18, 91, 27, -62, -3, 95, 35, 81, 108, 
        -108, 0, 52, -59, -36, -87, -64, 56, 48, 
        46, -60, -19, 2, 24, -71, 26, 43, 47, 
        -65, 58, 24, -39, 53, 49, 34, -5, 65, 
        -96, -41, 6, -85, -12, 84, -58, 36, 19, 
        -34, 86, -39, -1, -38, 73, -101, -87, 21, 
        42, 38, -13, -100, -88, 74, 53, -52, -93, 
        25, -70, -22, -94, 56, -15, 28, -122, -92, 
        -34, -76, -103, -29, -40, -18, 43, 18, -32, 
        -37, -85, 69, 15, 100, 38, -94, -50, -85, 
        73, 1, -60, 19, 80, 12, -68, -5, 60, 
        -89, -127, 65, -97, -33, -41, -6, -27, -126, 
        -59, 0, -26, -4, -23, -97, 59, -37, -44, 
        -81, -46, 69, -47, 5, 54, -29, -30, 106, 
        56, 59, -73, 104, 47, 94, 16, -83, 32, 
        93, 42, 79, 85, -15, -25, 5, 57, -95, 
        8, -52, -37, 73, 64, -45, 25, -70, 54, 
        -23, 38, -95, -121, 44, 61, -29, -81, 84, 
        -14, -56, -66, -109, 28, -46, -89, -37, 49, 
        -62, 57, -34, 33, -18, -124, -17, 1, -81, 
        -11, -18, -101, -52, 50, -54, -36, 6, 33, 
        -37, 8, -71, 83, -82, 9, 105, 66, -108, 
        52, -118, -89, -70, -37, -10, -105, 73, -103, 
        -77, -33, 54, 41, -31, -57, 94, 25, -89, 
        18, 32, 64, 45, 108, -34, 10, 98, 101, 
        54, 0, 50, 65, -22, 32, 27, -90, -56, 
        -51, 39, -77, -7, 34, 20, 59, -84, -2, 
        -111, 23, -87, -122, 56, 41, -85, -37, 76, 
        -31, 11, -28, -36, -12, -1, 5, -40, 7, 
        -19, 24, 28, -6, 0, -3, -60, -3, 37, 
        14, -13, 69, 28, -26, -5, -2, 0, -81, 
        28, 31, 1, -26, -5, 15, -9, 17, 2, 
        -8, 13, 18, -12, 20, 0, 10, -4, 14, 
        -5, -35, -60, -18, -24, -108, -22, -6, -92, 
        -38, -47, -34, 35, -16, -24, -18, 6, -64, 
        -16, 17, 14, 28, 16, -1, -27, -25, -23, 
        12, -24, 43, 4, -10, 0, 29, 14, -11, 
        11, 33, -10, -8, 1, 13, -28, 20, 13, 
        -26, -23, -26, 0, -8, 21, -26, -18, 13, 
        -7, -4, -21, -21, 42, 21, -42, -33, 33, 
        -8, -32, 6, 41, -64, 23, 54, -26, -38, 
        16, 2, -30, -16, -5, -13, 15, 10, 2, 
        -18, -11, -23, 3, 5, -33, -54, -8, 36, 
        17, 15, 22, -22, -2, 4, -60, -30, 28, 
        14, 35, 28, -35, -23, 9, -50, 20, 42, 
        77, -44, 69, 54, 52, -73, 64, -48, -127, 
        -30, 13, 9, -30, 4, -11, 25, 12, 29, 
        -10, 21, -29, 7, -11, -2, 18, 26, 16, 
        -6, 14, 17, -42, 9, -43, -25, -53, 6, 
        14, 50, 25, 11, 19, -47, 7, 51, 35, 
        -11, 31, 30, -37, 19, 61, -24, -58, 40, 
        -25, -10, -14, -32, 10, -14, -23, -18, -5, 
        -26, 32, 6, -18, 32, 1, -52, -37, 29, 
        3, -29, 4, -27, -8, 20, 17, 12, 4, 
        26, 91, 50, -37, 86, 101, -37, 13, 127, 
        -16, 1, 32, 24, -14, 9, -24, -25, -1, 
        9, -8, -18, 4, -19, -3, 27, -24, -18, 
        63, -21, -20, -10, -11, -46, 6, 55, 37, 
        37, 32, 107, 9, -19, 38, -39, -57, -9, 
        52, 33, -12, -10, 17, -21, 11, 62, 59
        }; 

        for (i = 0; i < (3 * 3 * 32 * 32 + 2); i = i + 4) begin
            ram.mem[1500 + (i / 4)][ 7: 0] = filter_data[8*((3 * 3 * 3 * 6 + 2) - 1 - i) +: 8];
            ram.mem[1500 + (i / 4)][15: 8] = filter_data[8*((3 * 3 * 3 * 6 + 2) - 2 - i) +: 8];
            ram.mem[1500 + (i / 4)][23:16] = filter_data[8*((3 * 3 * 3 * 6 + 2) - 3 - i) +: 8];
            ram.mem[1500 + (i / 4)][31:24] = filter_data[8*((3 * 3 * 3 * 6 + 2) - 4 - i) +: 8];
        end

        // Bias
        bias_data = {
            -28517, 2966, 5775, 5654, -11145, 7002, 8439, -9378, 8529, -489, -38044, -34300, 4925, -28784, -1970, 60, -8178, -26840, -28935, -31502, -10251, 6148, -3370, -8798, 7343, -44597, -6740, -31376, -15323, 3003, -31031, -2781
        };
        for (i = 0; i < BIS_SIZE; i = i + 1) begin
            ram.mem[1400 + i] = bias_data[32*(BIS_SIZE - 1 - i) +: 32];
        end

    end

`elsif CL_TC7
/* Test case 7 */
     /* 
        Description:
           - Input Feature Map's size : 13 x 13 x 32     => 5408
           - Kernel's size            : 3 x 3 x 32 x 3 => 9216
           - Output Feature Map's size: 11 x 11 x 3     => 150
           - Bias's size              : 3         =>  3872
           - Partial-Sum's size       : 6 x 6 x 6 x 4 => 864
    */

    localparam 
        IFM_SIZE = 28 * 28 * 3,
        KER_SIZE = 3 * 3 * 3 * 32,
        OFM_SIZE = 26 * 26 * 3,
        BIS_SIZE = 3,
        PAS_SIZE = 5 * 5 * 6;

    initial begin
        // al_accel_mem_read_ready = 1'b 0;
        // al_accel_mem_write_ready = 1'b 0;
        // #10
        // repeat (2000) @(posedge clk) begin
        //     #2 al_accel_mem_read_ready = $random;
        // end
        // #10 
        al_accel_mem_read_ready    = 1'b 1;
        al_accel_mem_write_ready   = 1'b 1;
    end

    initial begin
        al_accel_cfgreg_di   = 32'd 0; al_accel_cfgreg_sel = 5'd 0; 
        al_accel_cfgreg_wenb =  1'd 0;
        al_accel_flow_enb    =  1'b 0;
        #42
        al_accel_cfgreg_wenb =  1'd 1;
    // Config Data
        #10 // i_base_addr
        al_accel_cfgreg_di   = 32'd 0000;       al_accel_cfgreg_sel = 5'd 0; 

        #10 // kw_base_addr
        al_accel_cfgreg_di   = 32'd 6000;       al_accel_cfgreg_sel = 5'd 1; 

        #10 // o_base_addr
        al_accel_cfgreg_di   = 32'd 16000;       al_accel_cfgreg_sel = 5'd 2; 

        #10 // b_base_addr
        al_accel_cfgreg_di   = 32'd 5600;       al_accel_cfgreg_sel = 5'd 3; 

        #10 // ps_base_addr
        al_accel_cfgreg_di   = 32'd 20000;       al_accel_cfgreg_sel = 5'd 4; 

        #10 // {stride_height, stride_width, cfg_act_func_typ, cfg_layer_typ}
        al_accel_cfgreg_di   = {16'd 0, 4'd 1, 4'd 1, RELU, CONV}; al_accel_cfgreg_sel = 5'd 5; 

        #10 // {weight_kernel_patch_height, weight_kernel_patch_width}
        al_accel_cfgreg_di   = {16'd 3, 16'd 3}; al_accel_cfgreg_sel = 5'd 6; 

        #10 // {nok_ofm_depth, kernel_ifm_depth} 
        al_accel_cfgreg_di   = {16'd 3, 16'd 3}; al_accel_cfgreg_sel = 5'd 7;
        
        #10 // {ifm_height, ifm_width}  
        al_accel_cfgreg_di   = {16'd 28, 16'd 28}; al_accel_cfgreg_sel = 5'd 8;

        #10 // {ofm_height, ofm_width}
        al_accel_cfgreg_di   = {16'd 26, 16'd 26}; al_accel_cfgreg_sel = 5'd 9;

        #10 // {output2D_size, input2D_size}  
        al_accel_cfgreg_di   = {16'd 676, 16'd 784}; al_accel_cfgreg_sel = 5'd 10;

        #10 // kernel3D_size
        al_accel_cfgreg_di   = {16'd  0, 16'd 3}; al_accel_cfgreg_sel = 5'd 11;

        // Output Quantize Buffer
        #10 // output_quant_sel 0
        al_accel_cfgreg_di   = {24'd 0, 8'd 0} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2006707479 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 1
        al_accel_cfgreg_di   = {24'd 0, 8'd 1} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1433835724 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 2
        al_accel_cfgreg_di   = {24'd 0, 8'd 2} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1192390444 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 3
        al_accel_cfgreg_di   = {24'd 0, 8'd 3} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1361289408 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 4
        al_accel_cfgreg_di   = {24'd 0, 8'd 4} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1285031363 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 5
        al_accel_cfgreg_di   = {24'd 0, 8'd 5} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2063009507 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 6
        al_accel_cfgreg_di   = {24'd 0, 8'd 6} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2143833947 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 7
        al_accel_cfgreg_di   = {24'd 0, 8'd 7} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2040046477 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 11} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 8
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1117137979 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 9
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1529727281 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 10
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1118076866 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 11
        al_accel_cfgreg_di   = {24'd 0, 8'd 11} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1909265169 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 12
        al_accel_cfgreg_di   = {24'd 0, 8'd 12} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1213134709 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 13
        al_accel_cfgreg_di   = {24'd 0, 8'd 13} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1219315125 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 14
        al_accel_cfgreg_di   = {24'd 0, 8'd 14} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1693522756 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 15
        al_accel_cfgreg_di   = {24'd 0, 8'd 15} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1244537046 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 16
        al_accel_cfgreg_di   = {24'd 0, 8'd 16} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1439731708 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 17
        al_accel_cfgreg_di   = {24'd 0, 8'd 17} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1469553438 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 18
        al_accel_cfgreg_di   = {24'd 0, 8'd 18} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1858048416 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 11} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 19
        al_accel_cfgreg_di   = {24'd 0, 8'd 19} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1955939902 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 11} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 20
        al_accel_cfgreg_di   = {24'd 0, 8'd 20} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1424595433 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 21
        al_accel_cfgreg_di   = {24'd 0, 8'd 21} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1295986055 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 22
        al_accel_cfgreg_di   = {24'd 0, 8'd 22} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1959811992 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 23
        al_accel_cfgreg_di   = {24'd 0, 8'd 23} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1607690141 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 24
        al_accel_cfgreg_di   = {24'd 0, 8'd 24} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1265787593 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 25
        al_accel_cfgreg_di   = {24'd 0, 8'd 25} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1154422605 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 26
        al_accel_cfgreg_di   = {24'd 0, 8'd 26} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1891572973 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 27
        al_accel_cfgreg_di   = {24'd 0, 8'd 27} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1267784783 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 28
        al_accel_cfgreg_di   = {24'd 0, 8'd 28} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1192481101 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 10} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 29
        al_accel_cfgreg_di   = {24'd 0, 8'd 29} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1139166983 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 30
        al_accel_cfgreg_di   = {24'd 0, 8'd 30} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 1242432765 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 8} ; al_accel_cfgreg_sel = 5'd 14;

        #10 // output_quant_sel 31
        al_accel_cfgreg_di   = {24'd 0, 8'd 31} ; al_accel_cfgreg_sel = 5'd 12;
        #10 // output_multiplier
        al_accel_cfgreg_di   = 32'd 2027832722 ; al_accel_cfgreg_sel = 5'd 13;
        #10 // output_shift
        al_accel_cfgreg_di   = {24'd 0, 8'd 9} ; al_accel_cfgreg_sel = 5'd 14;

    // Data Offset
        #10 // {ofm_pool_height,  ofm_pool_width}
        al_accel_cfgreg_di   = {16'd 0, 16'd 0}; al_accel_cfgreg_sel = 5'd 15;
        #10 // output2D_pool_size
        al_accel_cfgreg_di   = 32'd 0; al_accel_cfgreg_sel = 5'd 16;

    // Flow Run
        #10
        al_accel_cfgreg_wenb =  1'd 0;
        #10 
        al_accel_flow_enb    =  1'd 1;
        // #1000
        // al_accel_flow_enb    =  1'd 0;
        // #200
        al_accel_flow_enb    =  1'd 1;
		// repeat (2000) @(posedge clk) begin
        //     #2 al_accel_flow_enb = $random;
        // end
        // #10 
        al_accel_flow_enb    =  1'd 1;
    end

    reg [IFM_SIZE    * 8 - 1:0] input_data ; // Size: 7 x 7 x 3
    reg [KER_SIZE * 8 - 1:0] filter_data; // Size: 3 x 3 x 3 x 6
    reg [ BIS_SIZE  *32              - 1:0] bias_data  ; // Size: 6
    integer i;
    initial begin
        for (i = 0; i < 32768; i = i + 1)
            ram.mem[i] = 32'd 0;

        // Input Initilization
        input_data = {
            /* z = 0 */
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd44, 8'd56, 8'd30, 8'd22, -8'd68, -8'd92, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd93, 8'd125, 8'd125, 8'd125, 8'd125, 8'd112, 8'd69, 8'd69, 8'd69, 8'd69, 8'd69, 8'd69, 8'd69, 8'd69, 8'd41, -8'd76, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd61, -8'd14, -8'd56, -8'd14, 8'd34, 8'd98, 8'd125, 8'd96, 8'd125, 8'd125, 8'd125, 8'd121, 8'd100, 8'd125, 8'd125, 8'd11, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd111, -8'd62, -8'd114, -8'd61, -8'd61, -8'd61, -8'd69, -8'd107, 8'd107, 8'd125, -8'd22, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd45, 8'd124, 8'd80, -8'd110, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd106, 8'd104, 8'd126, -8'd45, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd0, 8'd125, 8'd109, -8'd84, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd69, 8'd120, 8'd125, -8'd66, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd4, 8'd125, 8'd58, -8'd123, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd119, 8'd76, 8'd119, -8'd70, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd2, 8'd125, 8'd53, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd53, 8'd122, 8'd111, -8'd71, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd109, 8'd92, 8'd125, 8'd37, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd125, 8'd74, 8'd125, 8'd90, -8'd93, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd90, 8'd125, 8'd125, -8'd51, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd97, 8'd95, 8'd125, -8'd13, -8'd127, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 8'd4, 8'd125, 8'd125, -8'd76, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd67, 8'd113, 8'd125, 8'd125, -8'd76, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd7, 8'd125, 8'd125, 8'd90, -8'd88, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd7, 8'd125, 8'd78, -8'd110, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, 
            -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128, -8'd128,
        };


        for (i = 0; i < (28 * 28 * 3); i = i + 4) begin
            ram.mem[0 + (i / 4)][ 7: 0] = input_data[8*((28 * 28 * 3) - 1 - i) +: 8];
            ram.mem[0 + (i / 4)][15: 8] = input_data[8*((28 * 28 * 3) - 2 - i) +: 8];
            ram.mem[0 + (i / 4)][23:16] = input_data[8*((28 * 28 * 3) - 3 - i) +: 8];
            ram.mem[0 + (i / 4)][31:24] = input_data[8*((28 * 28 * 3) - 4 - i) +: 8];
        end
        

        // Kernel 
        filter_data = {
            /* channel 0 */
            -8'd72, -8'd127, -8'd17, 8'd90, 8'd41, 8'd67, 8'd102, 8'd103, 8'd67,
            8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0,
            8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0,

            /* channel 1 */
            8'd78, 8'd73, 8'd66, 8'd31, 8'd108, 8'd46, 8'd0, 8'd4, 8'd127,
            8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0,
            8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0,

            /* channel 2 */
            8'd93, 8'd15, -8'd83, 8'd68, -8'd26, -8'd102, 8'd24, -8'd127, -8'd85,
            8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0,
            8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0,

        };
 
        for (i = 0; i < (3 * 3 * 3 * 3 + 2); i = i + 4) begin
            ram.mem[1500 + (i / 4)][ 7: 0] = filter_data[8*((3 * 3 * 3 * 3 + 2) - 1 - i) +: 8];
            ram.mem[1500 + (i / 4)][15: 8] = filter_data[8*((3 * 3 * 3 * 3 + 2) - 2 - i) +: 8];
            ram.mem[1500 + (i / 4)][23:16] = filter_data[8*((3 * 3 * 3 * 3 + 2)- 3 - i) +: 8];
            ram.mem[1500 + (i / 4)][31:24] = filter_data[8*((3 * 3 * 3 * 3 + 2) - 4 - i) +: 8];
        end


        // Bias
        bias_data = {
            32'd32, -32'd959, 32'd13568
        };

        for (i = 0; i < 3; i = i + 1) begin
            ram.mem[1400 + i] = bias_data[32*(32 - 1 - i) +: 32];
        end
    end
/*******************/
`endif 

    // Module init
    al_accel uut (
        .al_accel_cfgreg_di     (al_accel_cfgreg_di),
        .al_accel_cfgreg_sel    (al_accel_cfgreg_sel),
        .al_accel_cfgreg_wenb   (al_accel_cfgreg_wenb),

        .al_accel_rdata         (al_accel_rdata),
        .al_accel_raddr         (al_accel_raddr),
        .al_accel_renb          (al_accel_renb),
        .al_accel_mem_read_ready    (al_accel_mem_read_ready),
        .al_accel_mem_write_ready   (al_accel_mem_write_ready),

        .al_accel_wdata         (al_accel_wdata),
        .al_accel_waddr         (al_accel_waddr),
        .al_accel_wenb          (al_accel_wenb),
        .al_accel_wstrb         (al_accel_wstrb),

        .al_accel_flow_enb      (al_accel_flow_enb),
        .al_accel_cal_fin       (al_accel_cal_fin),
        .al_accel_flow_resetn   (resetn),

        .clk    (clk),
        .resetn (resetn)
    );

    al_accel_mem ram (
        .renb   (al_accel_renb),
        .raddr  (al_accel_raddr[13:2]),
        .rdata  (al_accel_rdata),

        .wenb   (al_accel_wenb),
        .wstrb  (al_accel_wstrb),
        .waddr  (al_accel_waddr[13:2]),
        .wdata  (al_accel_wdata),

        .clk    (clk)
    );


    // Debug Info
    initial begin
        $dumpfile("accel_vcd/al_accel_tb.vcd");
        $dumpvars(0, al_accel_tb);

        repeat (`TIME_TO_REPEAT) begin
			repeat (2000) @(posedge clk);
		end
        // $display("FINISH LAYER");
        // for (i = 0; i < 4096; i = i + 1) begin
        //     $display("Addr %d [%d]: %d %d %d %d | %d | %h", i, (i << 2),
        //         $signed(ram.mem[i][ 7: 0]), 
        //         $signed(ram.mem[i][15: 8]), 
        //         $signed(ram.mem[i][23:16]), 
        //         $signed(ram.mem[i][31:24]),
        //         $signed(ram.mem[i]),
        //         $signed(ram.mem[i])
        //     ); 
        // end
        // $display("*************");
        $display("HARDWARE RESULT");
        for (i = 750; i < 750 + OFM_SIZE/4; i = i + 1) begin
            $display("%d %d %d %d", 
                $signed(ram.mem[i][ 7: 0]), 
                $signed(ram.mem[i][15: 8]), 
                $signed(ram.mem[i][23:16]), 
                $signed(ram.mem[i][31:24])
            ); 
        end
        $display("*************");
		$finish;
    end
endmodule

module al_accel_mem #(
	parameter integer WORDS = 8192
) (
    input              renb,
    input       [11:0] raddr,
    output reg  [31:0] rdata,

    input              wenb,
	input       [ 3:0] wstrb,
	input       [11:0] waddr,
	input       [31:0] wdata,
	
    input clk
);
	reg [31:0] mem [WORDS - 1:0];

	always @(posedge clk) begin
        if (renb)
            rdata <= mem[raddr];
        
        if (wenb) begin
            if (wstrb[0]) mem[waddr][ 7: 0] <= wdata[ 7: 0];
            if (wstrb[1]) mem[waddr][15: 8] <= wdata[15: 8];
            if (wstrb[2]) mem[waddr][23:16] <= wdata[23:16];
            if (wstrb[3]) mem[waddr][31:24] <= wdata[31:24];
        end
	end
endmodule

